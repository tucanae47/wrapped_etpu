* NGSPICE file created from wrapped_etpu.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt wrapped_etpu active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_100_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6914_ _6914_/A _3205_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__ebufn_8
XFILLER_70_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3988_ _3988_/A _3988_/B _3985_/Y vssd1 vssd1 vccd1 vccd1 _3989_/C sky130_fd_sc_hd__or3b_1
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6776_ _6532_/Q _6776_/D vssd1 vssd1 vccd1 vccd1 _6776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5727_ _6253_/A _5704_/X _5705_/X vssd1 vssd1 vccd1 vccd1 _5727_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5658_ _6685_/Q _5650_/X _5655_/X _5657_/X _5640_/X vssd1 vssd1 vccd1 vccd1 _6685_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4609_ _4620_/B _4609_/B vssd1 vssd1 vccd1 vccd1 _4611_/B sky130_fd_sc_hd__xor2_1
X_5589_ _5638_/A vssd1 vssd1 vccd1 vccd1 _5589_/X sky130_fd_sc_hd__clkbuf_2
X_6865__125 vssd1 vssd1 vccd1 vccd1 _6865__125/HI _6974_/A sky130_fd_sc_hd__conb_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4960_ _4960_/A vssd1 vssd1 vccd1 vccd1 _6537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4891_ _6512_/Q _4887_/X _4888_/X input39/X vssd1 vssd1 vccd1 vccd1 _6512_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3911_ _3941_/A _4257_/A _3908_/D _3910_/Y vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__a22o_1
X_6630_ _6799_/CLK _6630_/D vssd1 vssd1 vccd1 vccd1 _6630_/Q sky130_fd_sc_hd__dfxtp_1
X_3842_ _3855_/B _3842_/B vssd1 vssd1 vccd1 vccd1 _3843_/B sky130_fd_sc_hd__xnor2_1
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater71 _6799_/CLK vssd1 vssd1 vccd1 vccd1 _6795_/CLK sky130_fd_sc_hd__buf_12
X_6561_ _6562_/CLK _6561_/D vssd1 vssd1 vccd1 vccd1 _6899_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3773_ _3786_/B _3771_/Y _3750_/B _3750_/Y vssd1 vssd1 vccd1 vccd1 _3775_/B sky130_fd_sc_hd__o211a_1
X_5512_ _6672_/Q _5508_/X _5562_/S vssd1 vssd1 vccd1 vccd1 _5512_/X sky130_fd_sc_hd__mux2_1
X_6492_ _6795_/CLK _6492_/D vssd1 vssd1 vccd1 vccd1 _6492_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6849__109 vssd1 vssd1 vccd1 vccd1 _6849__109/HI _6958_/A sky130_fd_sc_hd__conb_1
XFILLER_105_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5443_ _5456_/A _5443_/B vssd1 vssd1 vccd1 vccd1 _5444_/A sky130_fd_sc_hd__and2_1
X_5374_ _5374_/A vssd1 vssd1 vccd1 vccd1 _5396_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4325_ _4325_/A _4325_/B _4350_/A vssd1 vssd1 vccd1 vccd1 _4326_/A sky130_fd_sc_hd__and3_1
X_6829__89 vssd1 vssd1 vccd1 vccd1 _6829__89/HI _6938_/A sky130_fd_sc_hd__conb_1
XFILLER_99_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4256_ _4252_/A _4254_/X _4255_/X vssd1 vssd1 vccd1 vccd1 _6373_/D sky130_fd_sc_hd__o21a_1
X_3207_ _3219_/A vssd1 vssd1 vccd1 vccd1 _3212_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4187_ _4187_/A _4187_/B vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__xnor2_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6759_ _6763_/CLK _6759_/D vssd1 vssd1 vccd1 vccd1 _6759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5090_ _6903_/A _5075_/X _5089_/X _5068_/X vssd1 vssd1 vccd1 vccd1 _6565_/D sky130_fd_sc_hd__o211a_1
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4070_/A _4072_/B _4069_/X vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__o21a_1
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4041_ _4042_/B _4042_/C _4042_/A vssd1 vssd1 vccd1 vccd1 _4043_/B sky130_fd_sc_hd__a21o_1
XFILLER_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5992_ _5969_/X _5990_/X _5991_/X vssd1 vssd1 vccd1 vccd1 _5992_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _5186_/A vssd1 vssd1 vccd1 vccd1 _5118_/B sky130_fd_sc_hd__buf_2
XFILLER_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6613_ _6667_/CLK _6613_/D vssd1 vssd1 vccd1 vccd1 _6613_/Q sky130_fd_sc_hd__dfxtp_1
X_4874_ _6500_/Q _4870_/X _4873_/X input36/X vssd1 vssd1 vccd1 vccd1 _6500_/D sky130_fd_sc_hd__a22o_1
X_3825_ _3847_/A _3825_/B vssd1 vssd1 vccd1 vccd1 _3825_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6544_ _6546_/CLK _6544_/D vssd1 vssd1 vccd1 vccd1 _6544_/Q sky130_fd_sc_hd__dfxtp_1
X_3756_ _3756_/A _3801_/A vssd1 vssd1 vccd1 vccd1 _3797_/A sky130_fd_sc_hd__or2_1
X_6475_ _6763_/CLK _6475_/D vssd1 vssd1 vccd1 vccd1 _6475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3687_ _3686_/A _3686_/B _3686_/C vssd1 vssd1 vccd1 vccd1 _3694_/C sky130_fd_sc_hd__a21o_1
X_5426_ _5439_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5427_/A sky130_fd_sc_hd__and2_1
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5357_ _6630_/Q _6629_/Q _5872_/A _6631_/Q _6632_/Q vssd1 vssd1 vccd1 vccd1 _5971_/B
+ sky130_fd_sc_hd__a2111oi_4
X_5288_ _6608_/Q _5294_/B vssd1 vssd1 vccd1 vccd1 _5289_/A sky130_fd_sc_hd__and2_1
X_4308_ _4517_/B vssd1 vssd1 vccd1 vccd1 _4479_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4239_ _4239_/A vssd1 vssd1 vccd1 vccd1 _4239_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ _4613_/A _4590_/B vssd1 vssd1 vccd1 vccd1 _4615_/D sky130_fd_sc_hd__xor2_1
X_3610_ _3759_/A _6653_/Q _3681_/D _3644_/D vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__and4_1
X_3541_ _3541_/A _3541_/B vssd1 vssd1 vccd1 vccd1 _3542_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3472_ _3472_/A vssd1 vssd1 vccd1 vccd1 _6314_/D sky130_fd_sc_hd__clkbuf_1
X_6260_ _6260_/A _6263_/B vssd1 vssd1 vccd1 vccd1 _6260_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5211_ _5044_/B _5210_/X _5088_/A vssd1 vssd1 vccd1 vccd1 _5212_/C sky130_fd_sc_hd__a21o_1
X_6191_ _6786_/Q _5342_/X _6188_/X _6190_/X vssd1 vssd1 vccd1 vccd1 _6786_/D sky130_fd_sc_hd__o211a_1
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5142_ _5142_/A vssd1 vssd1 vccd1 vccd1 _6574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5073_ _5047_/X _5071_/X _5072_/X _5055_/X vssd1 vssd1 vccd1 vccd1 _5073_/X sky130_fd_sc_hd__a31o_2
XFILLER_65_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4024_ _4024_/A _4024_/B vssd1 vssd1 vccd1 vccd1 _4024_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5975_ _6023_/A vssd1 vssd1 vccd1 vccd1 _6056_/B sky130_fd_sc_hd__clkbuf_2
X_4926_ _4925_/X _6530_/Q _4926_/S vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__mux2_1
X_4857_ _4857_/A vssd1 vssd1 vccd1 vccd1 _6490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3808_ _3836_/A _3835_/A _3808_/C _3808_/D vssd1 vssd1 vccd1 vccd1 _3809_/B sky130_fd_sc_hd__nand4_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6527_ _6528_/CLK _6527_/D vssd1 vssd1 vccd1 vccd1 _6527_/Q sky130_fd_sc_hd__dfxtp_1
X_4788_ _4788_/A vssd1 vssd1 vccd1 vccd1 _6459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3739_ _3703_/B _3703_/Y _3737_/Y _3738_/X vssd1 vssd1 vccd1 vccd1 _3741_/B sky130_fd_sc_hd__a211o_1
XFILLER_106_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6458_ _6789_/CLK _6458_/D vssd1 vssd1 vccd1 vccd1 _6458_/Q sky130_fd_sc_hd__dfxtp_1
X_6389_ _6795_/CLK _6389_/D vssd1 vssd1 vccd1 vccd1 _6389_/Q sky130_fd_sc_hd__dfxtp_1
X_5409_ _5406_/X _5707_/A _5409_/C vssd1 vssd1 vccd1 vccd1 _5410_/A sky130_fd_sc_hd__and3b_1
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5760_ _6701_/Q _5652_/X _5770_/S vssd1 vssd1 vccd1 vccd1 _5760_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ _6369_/Q _4711_/B vssd1 vssd1 vccd1 vccd1 _4712_/A sky130_fd_sc_hd__and2_1
X_5691_ _6688_/Q _3357_/X _5688_/X _5690_/X vssd1 vssd1 vccd1 vccd1 _6688_/D sky130_fd_sc_hd__o211a_1
X_4642_ _4642_/A _4642_/B _4642_/C vssd1 vssd1 vccd1 vccd1 _4644_/A sky130_fd_sc_hd__and3_1
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4573_ _4573_/A _4573_/B vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__nor2_2
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6312_ _6531_/CLK _6312_/D vssd1 vssd1 vccd1 vccd1 _6312_/Q sky130_fd_sc_hd__dfxtp_1
X_3524_ _3552_/A _5217_/D _3521_/D _3523_/Y vssd1 vssd1 vccd1 vccd1 _3524_/X sky130_fd_sc_hd__a22o_1
X_3455_ _3455_/A vssd1 vssd1 vccd1 vccd1 _6306_/D sky130_fd_sc_hd__clkbuf_1
X_6243_ _6243_/A _6243_/B vssd1 vssd1 vccd1 vccd1 _6243_/Y sky130_fd_sc_hd__nand2_1
X_3386_ _6292_/Q _6291_/Q _3385_/X _4259_/A vssd1 vssd1 vccd1 vccd1 _3392_/C sky130_fd_sc_hd__o31a_1
X_6174_ _6779_/Q _6169_/X _6173_/X _6165_/X vssd1 vssd1 vccd1 vccd1 _6779_/D sky130_fd_sc_hd__o211a_1
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5125_ _6910_/A _5149_/B vssd1 vssd1 vccd1 vccd1 _5129_/B sky130_fd_sc_hd__or2_1
XFILLER_84_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5056_ _5047_/X _5051_/X _5054_/X _5055_/X vssd1 vssd1 vccd1 vccd1 _5056_/X sky130_fd_sc_hd__a31o_1
X_4007_ _4036_/A _4057_/B _4036_/C vssd1 vssd1 vccd1 vccd1 _4009_/B sky130_fd_sc_hd__nand3_1
XFILLER_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5958_ _5935_/X _5956_/X _5957_/X _5687_/X vssd1 vssd1 vccd1 vccd1 _5958_/X sky130_fd_sc_hd__a211o_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _4919_/A _4909_/B vssd1 vssd1 vccd1 vccd1 _4909_/X sky130_fd_sc_hd__and2_1
XFILLER_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5889_ _5919_/A vssd1 vssd1 vccd1 vccd1 _5889_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_5 _3326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3243_/A vssd1 vssd1 vccd1 vccd1 _3240_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6930_ _6930_/A _3223_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6792_ _6799_/CLK _6792_/D vssd1 vssd1 vccd1 vccd1 _6792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5812_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5812_/X sky130_fd_sc_hd__clkbuf_2
X_5743_ _5915_/A vssd1 vssd1 vccd1 vccd1 _5743_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5674_ _6687_/Q _5650_/X _5671_/X _5673_/X _5640_/X vssd1 vssd1 vccd1 vccd1 _6687_/D
+ sky130_fd_sc_hd__o221a_1
X_4625_ _4637_/A _4636_/A _4636_/B _4637_/B vssd1 vssd1 vccd1 vccd1 _4626_/B sky130_fd_sc_hd__nand4_1
X_4556_ _4557_/A _4557_/B _4557_/C vssd1 vssd1 vccd1 vccd1 _4572_/A sky130_fd_sc_hd__o21ai_2
XFILLER_116_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3507_ _4259_/A vssd1 vssd1 vccd1 vccd1 _5162_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4487_ _4487_/A _4487_/B vssd1 vssd1 vccd1 vccd1 _4487_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3438_ _3792_/B vssd1 vssd1 vccd1 vccd1 _3808_/C sky130_fd_sc_hd__clkbuf_2
X_6226_ _6267_/A vssd1 vssd1 vccd1 vccd1 _6226_/X sky130_fd_sc_hd__clkbuf_2
X_3369_ _3375_/A _3368_/Y _6499_/D vssd1 vssd1 vccd1 vccd1 _6494_/D sky130_fd_sc_hd__o21a_1
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6157_ _6182_/B vssd1 vssd1 vccd1 vccd1 _6167_/B sky130_fd_sc_hd__clkbuf_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5108_/A _5108_/B vssd1 vssd1 vccd1 vccd1 _5108_/X sky130_fd_sc_hd__or2_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6088_ _6466_/Q _6081_/X _6070_/X _6087_/X _6482_/Q vssd1 vssd1 vccd1 vccd1 _6088_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_122_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5039_ _5011_/X _5037_/X _5038_/X _5019_/X vssd1 vssd1 vccd1 vccd1 _5039_/X sky130_fd_sc_hd__a31o_1
XFILLER_82_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4410_ _4410_/A _4426_/A vssd1 vssd1 vccd1 vccd1 _4411_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5390_ _5797_/A _5724_/S _6637_/Q vssd1 vssd1 vccd1 vccd1 _5391_/B sky130_fd_sc_hd__a21oi_1
XFILLER_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4341_ _4342_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__nand2_1
X_4272_ _4679_/A vssd1 vssd1 vccd1 vccd1 _4655_/B sky130_fd_sc_hd__clkbuf_4
X_3223_ _3224_/A vssd1 vssd1 vccd1 vccd1 _3223_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6011_ _6011_/A vssd1 vssd1 vccd1 vccd1 _6011_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6913_ _6913_/A _3204_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__ebufn_8
XFILLER_82_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3987_ _5193_/A vssd1 vssd1 vccd1 vccd1 _5239_/B sky130_fd_sc_hd__buf_4
X_6775_ _6532_/Q _6775_/D vssd1 vssd1 vccd1 vccd1 _6775_/Q sky130_fd_sc_hd__dfxtp_1
X_5726_ _5581_/X _5698_/X _5699_/X _5725_/X vssd1 vssd1 vccd1 vccd1 _5726_/X sky130_fd_sc_hd__o211a_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5657_ _6280_/A _5638_/X _5627_/X _5616_/X vssd1 vssd1 vccd1 vccd1 _5657_/X sky130_fd_sc_hd__a31o_1
X_4608_ _4588_/A _4588_/B _4607_/Y vssd1 vssd1 vccd1 vccd1 _4609_/B sky130_fd_sc_hd__a21boi_1
X_5588_ _6484_/Q vssd1 vssd1 vccd1 vccd1 _6253_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4539_ _4536_/X _4537_/X _4538_/Y vssd1 vssd1 vccd1 vccd1 _6391_/D sky130_fd_sc_hd__a21oi_1
XFILLER_89_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6209_ _6263_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6209_/X sky130_fd_sc_hd__or2_1
XFILLER_85_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4890_ _6511_/Q _4887_/X _4888_/X input38/X vssd1 vssd1 vccd1 vccd1 _6511_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3910_ _3928_/A vssd1 vssd1 vccd1 vccd1 _3910_/Y sky130_fd_sc_hd__inv_2
X_3841_ _3851_/A _3855_/A vssd1 vssd1 vccd1 vccd1 _3842_/B sky130_fd_sc_hd__nor2_1
Xrepeater72 _6799_/CLK vssd1 vssd1 vccd1 vccd1 _6667_/CLK sky130_fd_sc_hd__buf_12
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3772_ _3750_/B _3750_/Y _3786_/B _3771_/Y vssd1 vssd1 vccd1 vccd1 _3826_/A sky130_fd_sc_hd__a211oi_4
X_6560_ _6562_/CLK _6560_/D vssd1 vssd1 vccd1 vccd1 _6898_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5511_ _5669_/S vssd1 vssd1 vccd1 vccd1 _5562_/S sky130_fd_sc_hd__buf_2
X_6491_ _6795_/CLK _6491_/D vssd1 vssd1 vccd1 vccd1 _6491_/Q sky130_fd_sc_hd__dfxtp_2
X_6888__148 vssd1 vssd1 vccd1 vccd1 _6888__148/HI _6997_/A sky130_fd_sc_hd__conb_1
X_5442_ _3881_/A _3850_/A _5448_/S vssd1 vssd1 vccd1 vccd1 _5443_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5373_ _5373_/A vssd1 vssd1 vccd1 vccd1 _6633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4324_ _4324_/A _4324_/B vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__or2_2
XFILLER_99_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4255_ _5422_/A vssd1 vssd1 vccd1 vccd1 _4255_/X sky130_fd_sc_hd__buf_6
X_3206_ _3206_/A vssd1 vssd1 vccd1 vccd1 _3206_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4186_ _4207_/B _4186_/B vssd1 vssd1 vccd1 vccd1 _4187_/B sky130_fd_sc_hd__xnor2_4
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6758_ _6763_/CLK _6758_/D vssd1 vssd1 vccd1 vccd1 _6758_/Q sky130_fd_sc_hd__dfxtp_1
X_6689_ _6789_/CLK _6689_/D vssd1 vssd1 vccd1 vccd1 _6689_/Q sky130_fd_sc_hd__dfxtp_2
X_5709_ _6691_/Q _5553_/X _5764_/S vssd1 vssd1 vccd1 vccd1 _5709_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6580_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_4040_ _6661_/Q _4114_/C vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__and2_1
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5991_ _6481_/Q _6056_/B _5986_/X _5976_/X vssd1 vssd1 vccd1 vccd1 _5991_/X sky130_fd_sc_hd__a31o_1
XFILLER_92_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _5017_/A _5017_/B _5017_/C vssd1 vssd1 vccd1 vccd1 _5186_/A sky130_fd_sc_hd__and3_1
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6612_ _6667_/CLK _6612_/D vssd1 vssd1 vccd1 vccd1 _6612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4873_ _4873_/A vssd1 vssd1 vccd1 vccd1 _4873_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3824_ _3824_/A _3824_/B vssd1 vssd1 vccd1 vccd1 _3825_/B sky130_fd_sc_hd__nand2_1
X_6543_ _6584_/CLK _6543_/D vssd1 vssd1 vccd1 vccd1 _6543_/Q sky130_fd_sc_hd__dfxtp_1
X_3755_ _3787_/A _3755_/B _3755_/C _3755_/D vssd1 vssd1 vccd1 vccd1 _3801_/A sky130_fd_sc_hd__and4_1
XFILLER_118_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6474_ _6763_/CLK _6474_/D vssd1 vssd1 vccd1 vccd1 _6474_/Q sky130_fd_sc_hd__dfxtp_1
X_3686_ _3686_/A _3686_/B _3686_/C vssd1 vssd1 vccd1 vccd1 _3694_/B sky130_fd_sc_hd__nand3_1
XFILLER_118_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5425_ _5217_/B _3552_/A _5431_/S vssd1 vssd1 vccd1 vccd1 _5426_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5356_ _6647_/Q _3349_/X _6645_/Q _5882_/B vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__o31ai_4
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5287_ _5287_/A vssd1 vssd1 vccd1 vccd1 _6607_/D sky130_fd_sc_hd__clkbuf_1
X_4307_ _6667_/Q vssd1 vssd1 vccd1 vccd1 _4517_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4238_ _4219_/X _4220_/X _4235_/Y _4217_/Y vssd1 vssd1 vccd1 vccd1 _4238_/X sky130_fd_sc_hd__a211o_1
XFILLER_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4169_ _4169_/A _4169_/B _4169_/C vssd1 vssd1 vccd1 vccd1 _4169_/X sky130_fd_sc_hd__and3_1
XFILLER_83_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3540_ _3541_/A _3541_/B vssd1 vssd1 vccd1 vccd1 _3565_/A sky130_fd_sc_hd__or2_1
X_3471_ _6314_/Q _6518_/Q _3473_/S vssd1 vssd1 vccd1 vccd1 _3472_/A sky130_fd_sc_hd__mux2_1
X_5210_ _6703_/Q _6735_/Q _6767_/Q _6799_/Q _5188_/X _5014_/X vssd1 vssd1 vccd1 vccd1
+ _5210_/X sky130_fd_sc_hd__mux4_1
X_6190_ _6255_/A vssd1 vssd1 vccd1 vccd1 _6190_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5141_ _5160_/A _5141_/B _5141_/C vssd1 vssd1 vccd1 vccd1 _5142_/A sky130_fd_sc_hd__and3_1
X_5072_ _6808_/Q _5078_/B vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__or2_1
X_4023_ _4022_/B _4022_/C _4022_/A vssd1 vssd1 vccd1 vccd1 _4026_/B sky130_fd_sc_hd__o21ai_1
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _6736_/Q _5506_/X _5990_/S vssd1 vssd1 vccd1 vccd1 _5974_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4925_ _4928_/A _4925_/B vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__and2_1
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4856_ _6442_/Q _4856_/B vssd1 vssd1 vccd1 vccd1 _4857_/A sky130_fd_sc_hd__and2_1
X_3807_ _3835_/A _3808_/C _3808_/D _3836_/A vssd1 vssd1 vccd1 vccd1 _3809_/A sky130_fd_sc_hd__a22o_1
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6526_ _6528_/CLK _6526_/D vssd1 vssd1 vccd1 vccd1 _6526_/Q sky130_fd_sc_hd__dfxtp_1
X_4787_ _6411_/Q _4789_/B vssd1 vssd1 vccd1 vccd1 _4788_/A sky130_fd_sc_hd__and2_1
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3738_ _3750_/A _3750_/B _3750_/C vssd1 vssd1 vccd1 vccd1 _3738_/X sky130_fd_sc_hd__and3_1
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6457_ _6789_/CLK _6457_/D vssd1 vssd1 vccd1 vccd1 _6457_/Q sky130_fd_sc_hd__dfxtp_1
X_3669_ _3638_/X _3639_/X _3667_/X _3668_/Y vssd1 vssd1 vccd1 vccd1 _3669_/X sky130_fd_sc_hd__o211a_1
X_6388_ _6795_/CLK _6388_/D vssd1 vssd1 vccd1 vccd1 _6388_/Q sky130_fd_sc_hd__dfxtp_1
X_5408_ _5406_/B _5824_/A _5406_/A vssd1 vssd1 vccd1 vccd1 _5409_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5339_ _6222_/B vssd1 vssd1 vccd1 vccd1 _6192_/B sky130_fd_sc_hd__buf_2
XFILLER_87_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4710_/A vssd1 vssd1 vccd1 vccd1 _6424_/D sky130_fd_sc_hd__clkbuf_1
X_5690_ _5838_/A vssd1 vssd1 vccd1 vccd1 _5690_/X sky130_fd_sc_hd__clkbuf_2
X_4641_ _4641_/A vssd1 vssd1 vccd1 vccd1 _4642_/C sky130_fd_sc_hd__inv_2
XFILLER_30_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4572_ _4572_/A vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__inv_2
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6311_ _6531_/CLK _6311_/D vssd1 vssd1 vccd1 vccd1 _6311_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3523_ _3539_/A vssd1 vssd1 vccd1 vccd1 _3523_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3454_ _6306_/Q _6510_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _3455_/A sky130_fd_sc_hd__mux2_1
X_6242_ _6803_/Q _6226_/X _6241_/Y _6235_/X vssd1 vssd1 vccd1 vccd1 _6803_/D sky130_fd_sc_hd__o211a_1
X_3385_ _6294_/Q _6293_/Q _6295_/Q _3385_/D vssd1 vssd1 vccd1 vccd1 _3385_/X sky130_fd_sc_hd__or4_1
XFILLER_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6173_ _6273_/A _6180_/B vssd1 vssd1 vccd1 vccd1 _6173_/X sky130_fd_sc_hd__or2_1
X_5124_ _5186_/A vssd1 vssd1 vccd1 vccd1 _5149_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _5088_/A vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4006_ _4006_/A _4043_/A vssd1 vssd1 vccd1 vccd1 _4036_/C sky130_fd_sc_hd__nor2_1
XFILLER_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5957_ _6492_/Q _5957_/B _5957_/C vssd1 vssd1 vccd1 vccd1 _5957_/X sky130_fd_sc_hd__and3_1
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4908_ _4908_/A vssd1 vssd1 vccd1 vccd1 _6524_/D sky130_fd_sc_hd__clkbuf_1
X_5888_ _5946_/A vssd1 vssd1 vccd1 vccd1 _5888_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4839_ _6434_/Q _4845_/B vssd1 vssd1 vccd1 vccd1 _4840_/A sky130_fd_sc_hd__and2_1
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6509_ _6509_/CLK _6509_/D vssd1 vssd1 vccd1 vccd1 _6509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_6 _3330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5811_ _6708_/Q _5797_/X _5809_/X _5810_/X vssd1 vssd1 vccd1 vccd1 _6708_/D sky130_fd_sc_hd__o211a_1
X_6791_ _6809_/CLK _6791_/D vssd1 vssd1 vccd1 vccd1 _6791_/Q sky130_fd_sc_hd__dfxtp_1
X_5742_ _5610_/X _5741_/X _5757_/S vssd1 vssd1 vccd1 vccd1 _5742_/X sky130_fd_sc_hd__mux2_1
X_5673_ _6286_/A _5638_/X _6056_/C _5519_/X vssd1 vssd1 vccd1 vccd1 _5673_/X sky130_fd_sc_hd__a31o_1
X_4624_ _4637_/A _4636_/B _4597_/B _4636_/A vssd1 vssd1 vccd1 vccd1 _4626_/A sky130_fd_sc_hd__a22o_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4555_ _4584_/A _4555_/B vssd1 vssd1 vccd1 vccd1 _4557_/C sky130_fd_sc_hd__xnor2_2
X_3506_ _3506_/A vssd1 vssd1 vccd1 vccd1 _6334_/D sky130_fd_sc_hd__clkbuf_1
X_4486_ _4485_/A _4485_/B _4485_/C vssd1 vssd1 vccd1 vccd1 _4493_/C sky130_fd_sc_hd__a21o_1
X_6225_ _6264_/A vssd1 vssd1 vccd1 vccd1 _6267_/A sky130_fd_sc_hd__buf_2
X_3437_ _3755_/D vssd1 vssd1 vccd1 vccd1 _3792_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3368_ _6495_/Q _3370_/B _3405_/A vssd1 vssd1 vccd1 vccd1 _3368_/Y sky130_fd_sc_hd__nor3_1
XFILLER_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6156_ _6169_/A vssd1 vssd1 vccd1 vccd1 _6156_/X sky130_fd_sc_hd__clkbuf_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5107_ _6686_/Q _6718_/Q _6750_/Q _6782_/Q _5083_/X _4949_/A vssd1 vssd1 vccd1 vccd1
+ _5108_/B sky130_fd_sc_hd__mux4_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3299_ _3305_/A vssd1 vssd1 vccd1 vccd1 _3304_/A sky130_fd_sc_hd__buf_6
XFILLER_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6087_ _6113_/A vssd1 vssd1 vccd1 vccd1 _6087_/X sky130_fd_sc_hd__clkbuf_2
X_5038_ _6803_/Q _5044_/B vssd1 vssd1 vccd1 vccd1 _5038_/X sky130_fd_sc_hd__or2_1
XFILLER_26_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6989_ _6989_/A _3295_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4340_ _4340_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4342_/B sky130_fd_sc_hd__xnor2_1
XFILLER_113_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4271_ _4271_/A vssd1 vssd1 vccd1 vccd1 _6379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3222_ _3224_/A vssd1 vssd1 vccd1 vccd1 _3222_/Y sky130_fd_sc_hd__inv_2
X_6010_ _6742_/Q _5984_/X _6009_/X _5999_/X vssd1 vssd1 vccd1 vccd1 _6742_/D sky130_fd_sc_hd__o211a_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6912_ _6912_/A _3203_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__ebufn_8
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3986_ _3988_/A _3988_/B _3985_/Y vssd1 vssd1 vccd1 vccd1 _3986_/X sky130_fd_sc_hd__o21ba_1
X_6774_ _6532_/Q _6774_/D vssd1 vssd1 vccd1 vccd1 _6774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5725_ _5765_/A _5725_/B vssd1 vssd1 vccd1 vccd1 _5725_/X sky130_fd_sc_hd__or2_1
X_5656_ _6491_/Q vssd1 vssd1 vccd1 vccd1 _6280_/A sky130_fd_sc_hd__clkbuf_4
X_4607_ _4607_/A _4607_/B vssd1 vssd1 vccd1 vccd1 _4607_/Y sky130_fd_sc_hd__nand2_1
X_5587_ _5581_/X _5582_/X _5571_/X _5586_/X vssd1 vssd1 vccd1 vccd1 _5587_/X sky130_fd_sc_hd__o211a_1
XFILLER_116_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4538_ _4536_/X _4537_/X _3781_/X vssd1 vssd1 vccd1 vccd1 _4538_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4469_ _6671_/Q _6375_/Q _6376_/Q _6670_/Q vssd1 vssd1 vccd1 vccd1 _4473_/B sky130_fd_sc_hd__a22o_1
X_6208_ _6222_/B vssd1 vssd1 vccd1 vccd1 _6218_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6139_ _6767_/Q _6061_/X vssd1 vssd1 vccd1 vccd1 _6139_/X sky130_fd_sc_hd__or2b_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ _3840_/A _3840_/B vssd1 vssd1 vccd1 vccd1 _3855_/B sky130_fd_sc_hd__xnor2_2
X_3771_ _3785_/A _3769_/X _3728_/B _3751_/Y vssd1 vssd1 vccd1 vccd1 _3771_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5510_ _6637_/Q _6636_/Q _5510_/C vssd1 vssd1 vccd1 vccd1 _5669_/S sky130_fd_sc_hd__nor3_4
Xrepeater73 _6809_/CLK vssd1 vssd1 vccd1 vccd1 _6789_/CLK sky130_fd_sc_hd__buf_12
XFILLER_118_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6490_ _6795_/CLK _6490_/D vssd1 vssd1 vccd1 vccd1 _6490_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5441_ _5441_/A vssd1 vssd1 vccd1 vccd1 _5456_/A sky130_fd_sc_hd__clkbuf_2
X_5372_ _6633_/Q _5372_/B vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__and2_1
XFILLER_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4323_ _4324_/A _4324_/B vssd1 vssd1 vccd1 vccd1 _4325_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4254_ _4242_/A _4275_/A _4253_/X _4249_/A vssd1 vssd1 vccd1 vccd1 _4254_/X sky130_fd_sc_hd__a31o_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3205_ _3206_/A vssd1 vssd1 vccd1 vccd1 _3205_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4185_ _4155_/A _4154_/A _4154_/B vssd1 vssd1 vccd1 vccd1 _4186_/B sky130_fd_sc_hd__o21ba_2
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6871__131 vssd1 vssd1 vccd1 vccd1 _6871__131/HI _6980_/A sky130_fd_sc_hd__conb_1
XFILLER_23_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6757_ _6809_/CLK _6757_/D vssd1 vssd1 vccd1 vccd1 _6757_/Q sky130_fd_sc_hd__dfxtp_1
X_3969_ _4121_/B vssd1 vssd1 vccd1 vccd1 _4085_/B sky130_fd_sc_hd__clkbuf_2
X_5708_ _6690_/Q _5650_/X _5703_/X _5706_/X _5707_/X vssd1 vssd1 vccd1 vccd1 _6690_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6688_ _6789_/CLK _6688_/D vssd1 vssd1 vccd1 vccd1 _6688_/Q sky130_fd_sc_hd__dfxtp_2
X_5639_ _6273_/A _5638_/X _5627_/X _5616_/X vssd1 vssd1 vccd1 vccd1 _5639_/X sky130_fd_sc_hd__a31o_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6834__94 vssd1 vssd1 vccd1 vccd1 _6834__94/HI _6943_/A sky130_fd_sc_hd__conb_1
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5990_ _6739_/Q _5552_/X _5990_/S vssd1 vssd1 vccd1 vccd1 _5990_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4941_ _3324_/C _4962_/C _4941_/C _5008_/A vssd1 vssd1 vccd1 vccd1 _5017_/C sky130_fd_sc_hd__and4b_1
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4872_ _4895_/A vssd1 vssd1 vccd1 vccd1 _4873_/A sky130_fd_sc_hd__buf_2
X_6855__115 vssd1 vssd1 vccd1 vccd1 _6855__115/HI _6964_/A sky130_fd_sc_hd__conb_1
X_6611_ _6667_/CLK _6611_/D vssd1 vssd1 vccd1 vccd1 _6611_/Q sky130_fd_sc_hd__dfxtp_1
X_3823_ _3824_/A _3824_/B vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__or2_1
XFILLER_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6542_ _6551_/CLK _6542_/D vssd1 vssd1 vccd1 vccd1 _6542_/Q sky130_fd_sc_hd__dfxtp_1
X_3754_ _3755_/B _3755_/C _3792_/B _3787_/A vssd1 vssd1 vccd1 vccd1 _3756_/A sky130_fd_sc_hd__a22oi_1
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6473_ _6763_/CLK _6473_/D vssd1 vssd1 vccd1 vccd1 _6473_/Q sky130_fd_sc_hd__dfxtp_1
X_3685_ _3647_/A _3647_/B _3647_/C vssd1 vssd1 vccd1 vccd1 _3686_/C sky130_fd_sc_hd__a21bo_1
X_5424_ _5441_/A vssd1 vssd1 vccd1 vccd1 _5439_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5355_ _6635_/Q _6634_/Q _6633_/Q vssd1 vssd1 vccd1 vccd1 _5882_/B sky130_fd_sc_hd__nor3_2
X_5286_ _6607_/Q _5294_/B vssd1 vssd1 vccd1 vccd1 _5287_/A sky130_fd_sc_hd__and2_1
XFILLER_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4306_ _4306_/A vssd1 vssd1 vccd1 vccd1 _6384_/D sky130_fd_sc_hd__clkbuf_1
X_4237_ _4239_/A _4223_/B _4235_/Y _4236_/Y _3633_/X vssd1 vssd1 vccd1 vccd1 _6371_/D
+ sky130_fd_sc_hd__a311oi_1
XFILLER_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4168_ _4168_/A _4168_/B _4140_/A _4140_/B vssd1 vssd1 vccd1 vccd1 _4220_/C sky130_fd_sc_hd__or4bb_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4099_ _4074_/X _4062_/X _4097_/X _4098_/Y vssd1 vssd1 vccd1 vccd1 _4106_/B sky130_fd_sc_hd__o211ai_2
XFILLER_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6809_ _6809_/CLK _6809_/D vssd1 vssd1 vccd1 vccd1 _6809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3470_ _3470_/A vssd1 vssd1 vccd1 vccd1 _6313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5140_ _5119_/X _5139_/X _5115_/X vssd1 vssd1 vccd1 vccd1 _5141_/C sky130_fd_sc_hd__a21o_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5071_ _5077_/A _5071_/B vssd1 vssd1 vccd1 vccd1 _5071_/X sky130_fd_sc_hd__or2_1
XFILLER_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4022_ _4022_/A _4022_/B _4022_/C vssd1 vssd1 vccd1 vccd1 _4026_/A sky130_fd_sc_hd__or3_1
XFILLER_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5973_ _6048_/S vssd1 vssd1 vccd1 vccd1 _5990_/S sky130_fd_sc_hd__buf_2
X_4924_ _4924_/A vssd1 vssd1 vccd1 vccd1 _6529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4855_ _4855_/A vssd1 vssd1 vccd1 vccd1 _6489_/D sky130_fd_sc_hd__clkbuf_1
X_3806_ _3806_/A _3806_/B vssd1 vssd1 vccd1 vccd1 _3824_/A sky130_fd_sc_hd__or2_1
X_4786_ _4786_/A vssd1 vssd1 vccd1 vccd1 _6458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6525_ _6531_/CLK _6525_/D vssd1 vssd1 vccd1 vccd1 _6525_/Q sky130_fd_sc_hd__dfxtp_1
X_3737_ _3750_/B _3750_/C _3750_/A vssd1 vssd1 vccd1 vccd1 _3737_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6456_ _6789_/CLK _6456_/D vssd1 vssd1 vccd1 vccd1 _6456_/Q sky130_fd_sc_hd__dfxtp_1
X_3668_ _3664_/Y _3665_/X _3622_/B _3640_/Y vssd1 vssd1 vccd1 vccd1 _3668_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6387_ _6795_/CLK _6387_/D vssd1 vssd1 vccd1 vccd1 _6387_/Q sky130_fd_sc_hd__dfxtp_1
X_5407_ _5458_/A vssd1 vssd1 vccd1 vccd1 _5707_/A sky130_fd_sc_hd__buf_4
X_3599_ _3599_/A _3599_/B vssd1 vssd1 vccd1 vccd1 _3671_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5338_ _5870_/A _6143_/A vssd1 vssd1 vccd1 vccd1 _6222_/B sky130_fd_sc_hd__or2_1
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5269_ _6600_/Q _5271_/B vssd1 vssd1 vccd1 vccd1 _5270_/A sky130_fd_sc_hd__and2_1
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4640_ _4640_/A _4640_/B vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__xnor2_1
X_4571_ _4615_/B _4568_/X _4613_/B vssd1 vssd1 vccd1 vccd1 _4591_/A sky130_fd_sc_hd__o21bai_1
X_6310_ _6522_/CLK _6310_/D vssd1 vssd1 vccd1 vccd1 _6310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3522_ _3539_/B vssd1 vssd1 vccd1 vccd1 _3522_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3453_ _3499_/S vssd1 vssd1 vccd1 vccd1 _3462_/S sky130_fd_sc_hd__clkbuf_2
X_6241_ _6227_/X _6240_/Y _6230_/X vssd1 vssd1 vccd1 vccd1 _6241_/Y sky130_fd_sc_hd__o21ai_1
X_6172_ _6778_/Q _6169_/X _6171_/X _6165_/X vssd1 vssd1 vccd1 vccd1 _6778_/D sky130_fd_sc_hd__o211a_1
X_3384_ _6289_/Q _6290_/Q vssd1 vssd1 vccd1 vccd1 _3390_/C sky130_fd_sc_hd__and2_1
X_5123_ _5123_/A vssd1 vssd1 vccd1 vccd1 _6571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _6805_/Q _5078_/B vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__or2_1
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4005_ _4180_/B _6661_/Q _4039_/C _4005_/D vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__and4_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5956_ _5659_/X _5947_/X _5920_/A _5961_/B _6734_/Q vssd1 vssd1 vccd1 vccd1 _5956_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4907_ _4906_/X _6524_/Q _4910_/S vssd1 vssd1 vccd1 vccd1 _4908_/A sky130_fd_sc_hd__mux2_1
X_5887_ _6721_/Q _5850_/X _5886_/X _5863_/X vssd1 vssd1 vccd1 vccd1 _6721_/D sky130_fd_sc_hd__o211a_1
X_4838_ _4838_/A vssd1 vssd1 vccd1 vccd1 _6481_/D sky130_fd_sc_hd__clkbuf_1
X_4769_ _4791_/A vssd1 vssd1 vccd1 vccd1 _4778_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6508_ _6509_/CLK _6508_/D vssd1 vssd1 vccd1 vccd1 _6508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6439_ _6795_/CLK _6439_/D vssd1 vssd1 vccd1 vccd1 _6439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_7 _3330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6790_ _6809_/CLK _6790_/D vssd1 vssd1 vccd1 vccd1 _6790_/Q sky130_fd_sc_hd__dfxtp_1
X_5810_ _5838_/A vssd1 vssd1 vccd1 vccd1 _5810_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5741_ _6697_/Q _5611_/X _5751_/S vssd1 vssd1 vccd1 vccd1 _5741_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5672_ _6493_/Q vssd1 vssd1 vccd1 vccd1 _6286_/A sky130_fd_sc_hd__clkbuf_2
X_4623_ _4623_/A vssd1 vssd1 vccd1 vccd1 _4636_/A sky130_fd_sc_hd__clkbuf_2
X_4554_ _4554_/A _4585_/A vssd1 vssd1 vccd1 vccd1 _4555_/B sky130_fd_sc_hd__xnor2_1
X_3505_ _3639_/A _3865_/A _5008_/B vssd1 vssd1 vccd1 vccd1 _3506_/A sky130_fd_sc_hd__and3_1
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4485_ _4485_/A _4485_/B _4485_/C vssd1 vssd1 vccd1 vccd1 _4493_/B sky130_fd_sc_hd__nand3_2
X_6224_ _6224_/A _6224_/B _6224_/C vssd1 vssd1 vccd1 vccd1 _6264_/A sky130_fd_sc_hd__and3_2
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3436_ _6302_/Q vssd1 vssd1 vccd1 vccd1 _3755_/D sky130_fd_sc_hd__clkbuf_2
X_3367_ _6498_/Q _6497_/Q _6496_/Q vssd1 vssd1 vccd1 vccd1 _3405_/A sky130_fd_sc_hd__or3_1
X_6155_ _6772_/Q _6142_/X _6154_/X _6152_/X vssd1 vssd1 vccd1 vccd1 _6772_/D sky130_fd_sc_hd__o211a_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _6906_/A _5075_/X _5105_/X _5100_/X vssd1 vssd1 vccd1 vccd1 _6568_/D sky130_fd_sc_hd__o211a_1
XFILLER_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6086_ _6112_/A vssd1 vssd1 vccd1 vccd1 _6110_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3298_ _3298_/A vssd1 vssd1 vccd1 vccd1 _3298_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5037_ _5043_/A _5037_/B vssd1 vssd1 vccd1 vccd1 _5037_/X sky130_fd_sc_hd__or2_1
XFILLER_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6988_ _6988_/A _3294_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5939_ _5935_/X _5936_/X _5938_/X _5915_/X vssd1 vssd1 vccd1 vccd1 _5939_/X sky130_fd_sc_hd__a211o_1
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ _4270_/A _4270_/B vssd1 vssd1 vccd1 vccd1 _4271_/A sky130_fd_sc_hd__and2_1
XFILLER_113_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3221_ _3224_/A vssd1 vssd1 vccd1 vccd1 _3221_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6911_ _6911_/A _3202_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__ebufn_8
XFILLER_54_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6773_ _6809_/CLK _6773_/D vssd1 vssd1 vccd1 vccd1 _6773_/Q sky130_fd_sc_hd__dfxtp_1
X_3985_ _3985_/A _3985_/B vssd1 vssd1 vccd1 vccd1 _3985_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5724_ _6694_/Q _5584_/X _5724_/S vssd1 vssd1 vccd1 vccd1 _5725_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5655_ _5651_/X _5631_/X _5620_/X _5654_/X vssd1 vssd1 vccd1 vccd1 _5655_/X sky130_fd_sc_hd__o211a_1
X_4606_ _4606_/A _4642_/A vssd1 vssd1 vccd1 vccd1 _4620_/B sky130_fd_sc_hd__nor2_1
X_5586_ _5624_/A _5586_/B vssd1 vssd1 vccd1 vccd1 _5586_/X sky130_fd_sc_hd__or2_1
XFILLER_117_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4537_ _4505_/X _4615_/A _4566_/A vssd1 vssd1 vccd1 vccd1 _4537_/X sky130_fd_sc_hd__o21ba_1
X_4468_ _4468_/A _4468_/B _4468_/C vssd1 vssd1 vccd1 vccd1 _4468_/X sky130_fd_sc_hd__and3_1
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6207_ _6207_/A vssd1 vssd1 vccd1 vccd1 _6207_/X sky130_fd_sc_hd__clkbuf_2
X_3419_ _3419_/A vssd1 vssd1 vccd1 vccd1 _6298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4399_ _4623_/A _4373_/D _4400_/D _4547_/A vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__a22oi_1
X_6138_ _5667_/X _6493_/Q _6138_/S vssd1 vssd1 vccd1 vccd1 _6138_/X sky130_fd_sc_hd__mux2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _6096_/A vssd1 vssd1 vccd1 vccd1 _6070_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3770_ _3728_/B _3751_/Y _3785_/A _3769_/X vssd1 vssd1 vccd1 vccd1 _3786_/B sky130_fd_sc_hd__o211a_1
Xrepeater74 _6799_/CLK vssd1 vssd1 vccd1 vccd1 _6809_/CLK sky130_fd_sc_hd__buf_12
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5440_ _5440_/A vssd1 vssd1 vccd1 vccd1 _6654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5371_ _5371_/A vssd1 vssd1 vccd1 vccd1 _6632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4322_ _4296_/X _4304_/B _4320_/Y _4349_/A vssd1 vssd1 vccd1 vccd1 _4324_/B sky130_fd_sc_hd__o31ai_1
X_4253_ _4241_/A _4273_/A _4245_/B vssd1 vssd1 vccd1 vccd1 _4253_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3204_ _3206_/A vssd1 vssd1 vccd1 vccd1 _3204_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4184_ _4184_/A _4205_/B vssd1 vssd1 vccd1 vccd1 _4207_/B sky130_fd_sc_hd__nor2_2
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3968_ _6659_/Q vssd1 vssd1 vccd1 vccd1 _4121_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6756_ _6763_/CLK _6756_/D vssd1 vssd1 vccd1 vccd1 _6756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5707_ _5707_/A vssd1 vssd1 vccd1 vccd1 _5707_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6687_ _6799_/CLK _6687_/D vssd1 vssd1 vccd1 vccd1 _6687_/Q sky130_fd_sc_hd__dfxtp_1
X_3899_ _3899_/A _3899_/B _3913_/A vssd1 vssd1 vccd1 vccd1 _3900_/A sky130_fd_sc_hd__and3_1
X_5638_ _5638_/A vssd1 vssd1 vccd1 vccd1 _5638_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5569_ _6676_/Q _5551_/X _5564_/X _5568_/X _5540_/X vssd1 vssd1 vccd1 vccd1 _6676_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4940_ _6536_/Q _6331_/Q _5081_/A vssd1 vssd1 vccd1 vccd1 _4962_/C sky130_fd_sc_hd__and3b_1
X_4871_ _4929_/S _4867_/B vssd1 vssd1 vccd1 vccd1 _4895_/A sky130_fd_sc_hd__nor2b_4
X_6610_ _6667_/CLK _6610_/D vssd1 vssd1 vccd1 vccd1 _6610_/Q sky130_fd_sc_hd__dfxtp_1
X_3822_ _3833_/B _3822_/B vssd1 vssd1 vccd1 vccd1 _3824_/B sky130_fd_sc_hd__xor2_1
X_6541_ _6546_/CLK _6541_/D vssd1 vssd1 vccd1 vccd1 _6541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3753_ _3753_/A vssd1 vssd1 vccd1 vccd1 _3787_/A sky130_fd_sc_hd__clkbuf_2
X_6472_ _6763_/CLK _6472_/D vssd1 vssd1 vccd1 vccd1 _6472_/Q sky130_fd_sc_hd__dfxtp_1
X_3684_ _3684_/A _3684_/B _3684_/C vssd1 vssd1 vccd1 vccd1 _3686_/B sky130_fd_sc_hd__nand3_1
X_5423_ _5423_/A vssd1 vssd1 vccd1 vccd1 _6649_/D sky130_fd_sc_hd__clkbuf_1
X_5354_ _5824_/A vssd1 vssd1 vccd1 vccd1 _5797_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4305_ _4325_/A _4305_/B _4324_/A vssd1 vssd1 vccd1 vccd1 _4306_/A sky130_fd_sc_hd__and3_1
XFILLER_114_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5285_ _5374_/A vssd1 vssd1 vccd1 vccd1 _5294_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4236_ _4239_/A _4223_/B _4235_/Y vssd1 vssd1 vccd1 vccd1 _4236_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4167_ _4218_/B _4167_/B vssd1 vssd1 vccd1 vccd1 _4220_/B sky130_fd_sc_hd__or2_1
XFILLER_55_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4098_ _4098_/A _4098_/B _4098_/C vssd1 vssd1 vccd1 vccd1 _4098_/Y sky130_fd_sc_hd__nand3_2
XFILLER_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6808_ _6809_/CLK _6808_/D vssd1 vssd1 vccd1 vccd1 _6808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6739_ _6809_/CLK _6739_/D vssd1 vssd1 vccd1 vccd1 _6739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6878__138 vssd1 vssd1 vccd1 vccd1 _6878__138/HI _6987_/A sky130_fd_sc_hd__conb_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5070_ _6680_/Q _6712_/Q _6744_/Q _6776_/Q _5049_/X _5063_/X vssd1 vssd1 vccd1 vccd1
+ _5071_/B sky130_fd_sc_hd__mux4_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4021_ _4067_/B _4067_/C _4067_/A vssd1 vssd1 vccd1 vccd1 _4022_/C sky130_fd_sc_hd__o21a_1
XFILLER_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5972_ _5972_/A _6068_/A vssd1 vssd1 vccd1 vccd1 _6048_/S sky130_fd_sc_hd__nor2_2
X_4923_ _4922_/X _6529_/Q _4926_/S vssd1 vssd1 vccd1 vccd1 _4924_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4854_ _6441_/Q _4856_/B vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__and2_1
XFILLER_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3805_ _4990_/A _3805_/B vssd1 vssd1 vccd1 vccd1 _6345_/D sky130_fd_sc_hd__nor2_1
X_4785_ _6410_/Q _4789_/B vssd1 vssd1 vccd1 vccd1 _4786_/A sky130_fd_sc_hd__and2_1
X_6524_ _6531_/CLK _6524_/D vssd1 vssd1 vccd1 vccd1 _6524_/Q sky130_fd_sc_hd__dfxtp_1
X_3736_ _3552_/A _3808_/C _3692_/B _3691_/B vssd1 vssd1 vccd1 vccd1 _3750_/A sky130_fd_sc_hd__a31o_1
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3667_ _3667_/A vssd1 vssd1 vccd1 vccd1 _3667_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6455_ _6789_/CLK _6455_/D vssd1 vssd1 vccd1 vccd1 _6455_/Q sky130_fd_sc_hd__dfxtp_1
X_5406_ _5406_/A _5406_/B _5406_/C vssd1 vssd1 vccd1 vccd1 _5406_/X sky130_fd_sc_hd__and3_1
X_6386_ _6795_/CLK _6386_/D vssd1 vssd1 vccd1 vccd1 _6386_/Q sky130_fd_sc_hd__dfxtp_1
X_3598_ _3598_/A vssd1 vssd1 vccd1 vccd1 _3625_/A sky130_fd_sc_hd__inv_2
XFILLER_87_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5337_ _6268_/A _5337_/B vssd1 vssd1 vccd1 vccd1 _6143_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5268_ _5268_/A vssd1 vssd1 vccd1 vccd1 _6599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4219_ _4220_/B _4170_/Y _4220_/D _4218_/Y _4194_/B vssd1 vssd1 vccd1 vccd1 _4219_/X
+ sky130_fd_sc_hd__o32a_2
X_5199_ _6922_/A _5209_/B vssd1 vssd1 vccd1 vccd1 _5202_/B sky130_fd_sc_hd__or2_1
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4570_ _4615_/B _4568_/X _4569_/Y vssd1 vssd1 vccd1 vccd1 _6392_/D sky130_fd_sc_hd__a21oi_1
X_3521_ _3539_/A _5217_/D _3552_/A _3521_/D vssd1 vssd1 vccd1 vccd1 _3539_/B sky130_fd_sc_hd__and4b_1
XFILLER_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6240_ _6240_/A _6243_/B vssd1 vssd1 vccd1 vccd1 _6240_/Y sky130_fd_sc_hd__nand2_1
X_3452_ _3452_/A vssd1 vssd1 vccd1 vccd1 _6305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3383_ _3383_/A vssd1 vssd1 vccd1 vccd1 _6290_/D sky130_fd_sc_hd__clkbuf_1
X_6171_ _6270_/A _6180_/B vssd1 vssd1 vccd1 vccd1 _6171_/X sky130_fd_sc_hd__or2_1
XFILLER_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5122_ _5129_/A _5122_/B _5122_/C vssd1 vssd1 vccd1 vccd1 _5123_/A sky130_fd_sc_hd__and3_1
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _5181_/A vssd1 vssd1 vccd1 vccd1 _5078_/B sky130_fd_sc_hd__buf_2
XFILLER_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4004_ _6662_/Q vssd1 vssd1 vccd1 vccd1 _4180_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5955_ _6733_/Q _5946_/X _5954_/X _5933_/X vssd1 vssd1 vccd1 vccd1 _6733_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _4919_/A _4906_/B vssd1 vssd1 vccd1 vccd1 _4906_/X sky130_fd_sc_hd__and2_1
X_5886_ _6233_/A _5964_/D _5638_/A _5885_/X _5538_/X vssd1 vssd1 vccd1 vccd1 _5886_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4837_ _6433_/Q _4845_/B vssd1 vssd1 vccd1 vccd1 _4838_/A sky130_fd_sc_hd__and2_1
X_4768_ _4768_/A vssd1 vssd1 vccd1 vccd1 _6450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3719_ _3759_/A _3720_/C _3720_/D _6655_/Q vssd1 vssd1 vccd1 vccd1 _3722_/C sky130_fd_sc_hd__a22o_1
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6507_ _6509_/CLK _6507_/D vssd1 vssd1 vccd1 vccd1 _6507_/Q sky130_fd_sc_hd__dfxtp_1
X_4699_ _4699_/A vssd1 vssd1 vccd1 vccd1 _6419_/D sky130_fd_sc_hd__clkbuf_1
X_6438_ _6795_/CLK _6438_/D vssd1 vssd1 vccd1 vccd1 _6438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6369_ _6763_/CLK _6369_/D vssd1 vssd1 vccd1 vccd1 _6369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_8 _3330_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5740_ _6696_/Q _5718_/X _5738_/X _5739_/X vssd1 vssd1 vccd1 vccd1 _6696_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5667_/X _5631_/X _5620_/A _5670_/X vssd1 vssd1 vccd1 vccd1 _5671_/X sky130_fd_sc_hd__o211a_1
XFILLER_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4622_ _4622_/A vssd1 vssd1 vccd1 vccd1 _4637_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4553_ _4553_/A _4553_/B vssd1 vssd1 vccd1 vccd1 _4585_/A sky130_fd_sc_hd__and2_1
X_3504_ _5193_/A vssd1 vssd1 vccd1 vccd1 _5008_/B sky130_fd_sc_hd__clkbuf_8
X_4484_ _4445_/A _4445_/C _4445_/B vssd1 vssd1 vccd1 vccd1 _4485_/C sky130_fd_sc_hd__a21bo_1
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6223_ _6799_/Q _6207_/A _6222_/X _6216_/X vssd1 vssd1 vccd1 vccd1 _6799_/D sky130_fd_sc_hd__o211a_1
X_3435_ _3435_/A vssd1 vssd1 vccd1 vccd1 _6301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3366_ _6330_/Q _4993_/C _3340_/X vssd1 vssd1 vccd1 vccd1 _6332_/D sky130_fd_sc_hd__o21a_1
XFILLER_97_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6154_ _6243_/A _6154_/B vssd1 vssd1 vccd1 vccd1 _6154_/X sky130_fd_sc_hd__or2_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5105_ _5081_/X _5103_/X _5104_/X _5088_/X vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__a31o_1
XFILLER_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3297_ _3298_/A vssd1 vssd1 vccd1 vccd1 _3297_/Y sky130_fd_sc_hd__inv_2
X_6085_ _6085_/A vssd1 vssd1 vccd1 vccd1 _6755_/D sky130_fd_sc_hd__clkbuf_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _6675_/Q _6707_/Q _6739_/Q _6771_/Q _5012_/X _5029_/X vssd1 vssd1 vccd1 vccd1
+ _5037_/B sky130_fd_sc_hd__mux4_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6987_ _6987_/A _3292_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5938_ _6488_/Q _5957_/B _5943_/C vssd1 vssd1 vccd1 vccd1 _5938_/X sky130_fd_sc_hd__and3_1
XFILLER_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5869_ _6719_/Q _5850_/X _5868_/X _5863_/X vssd1 vssd1 vccd1 vccd1 _6719_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6570_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_3220_ _3224_/A vssd1 vssd1 vccd1 vccd1 _3220_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6910_ _6910_/A _3200_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__ebufn_8
XFILLER_82_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6772_ _6809_/CLK _6772_/D vssd1 vssd1 vccd1 vccd1 _6772_/Q sky130_fd_sc_hd__dfxtp_1
X_3984_ _4024_/A _4024_/B vssd1 vssd1 vccd1 vccd1 _3985_/B sky130_fd_sc_hd__xor2_1
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5723_ _6693_/Q _5718_/X _5722_/X _5690_/X vssd1 vssd1 vccd1 vccd1 _6693_/D sky130_fd_sc_hd__o211a_1
X_5654_ _5670_/A _5654_/B vssd1 vssd1 vccd1 vccd1 _5654_/X sky130_fd_sc_hd__or2_1
X_4605_ _4605_/A _4605_/B vssd1 vssd1 vccd1 vccd1 _4642_/A sky130_fd_sc_hd__nor2_1
X_5585_ _6678_/Q _5584_/X _5612_/S vssd1 vssd1 vccd1 vccd1 _5586_/B sky130_fd_sc_hd__mux2_1
X_4536_ _4566_/C _4566_/D vssd1 vssd1 vccd1 vccd1 _4536_/X sky130_fd_sc_hd__or2_1
XFILLER_117_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4467_ _4426_/X _4427_/X _4466_/A _4457_/X vssd1 vssd1 vccd1 vccd1 _4467_/X sky130_fd_sc_hd__a211o_1
X_4398_ _4576_/B vssd1 vssd1 vccd1 vccd1 _4623_/A sky130_fd_sc_hd__clkbuf_2
X_6206_ _6792_/Q _6194_/X _6205_/X _6203_/X vssd1 vssd1 vccd1 vccd1 _6792_/D sky130_fd_sc_hd__o211a_1
X_3418_ _5217_/B _6502_/Q _3427_/S vssd1 vssd1 vccd1 vccd1 _3419_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3349_ _6646_/Q vssd1 vssd1 vccd1 vccd1 _3349_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6137_ _6137_/A vssd1 vssd1 vccd1 vccd1 _6766_/D sky130_fd_sc_hd__clkbuf_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _6068_/A _6113_/A vssd1 vssd1 vccd1 vccd1 _6096_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5019_ _5088_/A vssd1 vssd1 vccd1 vccd1 _5019_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater75 _6532_/Q vssd1 vssd1 vccd1 vccd1 _6799_/CLK sky130_fd_sc_hd__buf_12
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5370_ _6632_/Q _5372_/B vssd1 vssd1 vccd1 vccd1 _5371_/A sky130_fd_sc_hd__and2_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4321_ _4296_/X _4304_/B _4320_/Y vssd1 vssd1 vccd1 vccd1 _4349_/A sky130_fd_sc_hd__o21ai_2
X_4252_ _4252_/A _4252_/B vssd1 vssd1 vccd1 vccd1 _6372_/D sky130_fd_sc_hd__nor2_1
X_3203_ _3206_/A vssd1 vssd1 vccd1 vccd1 _3203_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4183_ _4202_/A _4183_/B _4183_/C vssd1 vssd1 vccd1 vccd1 _4205_/B sky130_fd_sc_hd__and3_1
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6755_ _6809_/CLK _6755_/D vssd1 vssd1 vccd1 vccd1 _6755_/Q sky130_fd_sc_hd__dfxtp_1
X_3967_ _3967_/A _3967_/B vssd1 vssd1 vccd1 vccd1 _3995_/A sky130_fd_sc_hd__xnor2_1
X_5706_ _6237_/A _5704_/X _5705_/X vssd1 vssd1 vccd1 vccd1 _5706_/X sky130_fd_sc_hd__a21o_1
X_6686_ _6799_/CLK _6686_/D vssd1 vssd1 vccd1 vccd1 _6686_/Q sky130_fd_sc_hd__dfxtp_1
X_3898_ _3992_/A _4056_/A _4257_/A _4262_/A vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__nand4_2
X_5637_ _6489_/Q vssd1 vssd1 vccd1 vccd1 _6273_/A sky130_fd_sc_hd__clkbuf_4
X_5568_ _6243_/A _5534_/X _6286_/B _5567_/X vssd1 vssd1 vccd1 vccd1 _5568_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4519_ _4519_/A _6381_/Q vssd1 vssd1 vccd1 vccd1 _4541_/B sky130_fd_sc_hd__nand2_1
XFILLER_120_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5499_ _6622_/Q _5499_/B vssd1 vssd1 vccd1 vccd1 _5870_/B sky130_fd_sc_hd__or2_2
XFILLER_78_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4870_ _4870_/A vssd1 vssd1 vccd1 vccd1 _4870_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3821_ _3801_/A _3801_/B _3820_/Y vssd1 vssd1 vccd1 vccd1 _3822_/B sky130_fd_sc_hd__a21boi_1
X_6540_ _6546_/CLK _6540_/D vssd1 vssd1 vccd1 vccd1 _6540_/Q sky130_fd_sc_hd__dfxtp_1
X_3752_ _3769_/A _3752_/B _3730_/X vssd1 vssd1 vccd1 vccd1 _3769_/B sky130_fd_sc_hd__nor3b_1
X_6471_ _6763_/CLK _6471_/D vssd1 vssd1 vccd1 vccd1 _6471_/Q sky130_fd_sc_hd__dfxtp_1
X_3683_ _3684_/B _3684_/C _3684_/A vssd1 vssd1 vccd1 vccd1 _3686_/A sky130_fd_sc_hd__a21o_1
X_5422_ _5422_/A _5422_/B vssd1 vssd1 vccd1 vccd1 _5423_/A sky130_fd_sc_hd__and2_1
X_5353_ _6102_/A vssd1 vssd1 vccd1 vccd1 _5824_/A sky130_fd_sc_hd__buf_2
X_4304_ _4304_/A _4304_/B _4304_/C vssd1 vssd1 vccd1 vccd1 _4324_/A sky130_fd_sc_hd__or3_1
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5284_ _5284_/A vssd1 vssd1 vccd1 vccd1 _5374_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4235_ _4235_/A _4235_/B vssd1 vssd1 vccd1 vccd1 _4235_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4166_ _4218_/A _4164_/X _4135_/B _4169_/B vssd1 vssd1 vccd1 vccd1 _4167_/B sky130_fd_sc_hd__o211a_1
X_6825__85 vssd1 vssd1 vccd1 vccd1 _6825__85/HI _6934_/A sky130_fd_sc_hd__conb_1
XFILLER_83_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4097_ _4098_/B _4098_/C _4098_/A vssd1 vssd1 vccd1 vccd1 _4097_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6807_ _6809_/CLK _6807_/D vssd1 vssd1 vccd1 vccd1 _6807_/Q sky130_fd_sc_hd__dfxtp_1
X_4999_ _5129_/A _4999_/B _4999_/C vssd1 vssd1 vccd1 vccd1 _5000_/A sky130_fd_sc_hd__and3_1
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6738_ _6809_/CLK _6738_/D vssd1 vssd1 vccd1 vccd1 _6738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6669_ _6795_/CLK _6669_/D vssd1 vssd1 vccd1 vccd1 _6669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6861__121 vssd1 vssd1 vccd1 vccd1 _6861__121/HI _6970_/A sky130_fd_sc_hd__conb_1
XFILLER_96_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4020_ _4067_/A _4067_/B _4067_/C vssd1 vssd1 vccd1 vccd1 _4022_/B sky130_fd_sc_hd__nor3_1
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5971_ _5971_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _6068_/A sky130_fd_sc_hd__nand2_2
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4922_ _4928_/A _4922_/B vssd1 vssd1 vccd1 vccd1 _4922_/X sky130_fd_sc_hd__and2_1
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4853_ _4853_/A vssd1 vssd1 vccd1 vccd1 _6488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4784_ _4784_/A vssd1 vssd1 vccd1 vccd1 _6457_/D sky130_fd_sc_hd__clkbuf_1
X_3804_ _3804_/A _3828_/D vssd1 vssd1 vccd1 vccd1 _3805_/B sky130_fd_sc_hd__xor2_1
X_6523_ _6523_/CLK _6523_/D vssd1 vssd1 vccd1 vccd1 _6523_/Q sky130_fd_sc_hd__dfxtp_1
X_3735_ _3734_/A _3734_/B _3734_/C vssd1 vssd1 vccd1 vccd1 _3750_/C sky130_fd_sc_hd__a21o_1
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6454_ _6789_/CLK _6454_/D vssd1 vssd1 vccd1 vccd1 _6454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5405_ _5879_/A _5405_/B vssd1 vssd1 vccd1 vccd1 _6644_/D sky130_fd_sc_hd__nor2_1
X_3666_ _3622_/B _3640_/Y _3664_/Y _3665_/X vssd1 vssd1 vccd1 vccd1 _3667_/A sky130_fd_sc_hd__a211o_1
X_6385_ _6795_/CLK _6385_/D vssd1 vssd1 vccd1 vccd1 _6385_/Q sky130_fd_sc_hd__dfxtp_1
X_3597_ _3659_/A _3808_/D _3576_/A _3596_/X vssd1 vssd1 vccd1 vccd1 _3598_/A sky130_fd_sc_hd__a31o_1
X_5336_ _5876_/B _5880_/B vssd1 vssd1 vccd1 vccd1 _5870_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5267_ _6599_/Q _5271_/B vssd1 vssd1 vccd1 vccd1 _5268_/A sky130_fd_sc_hd__and2_1
XFILLER_102_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4218_ _4218_/A _4218_/B vssd1 vssd1 vccd1 vccd1 _4218_/Y sky130_fd_sc_hd__nor2_1
X_5198_ _5198_/A vssd1 vssd1 vccd1 vccd1 _6583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4149_ _4177_/A _4149_/B _4183_/B _6357_/Q vssd1 vssd1 vccd1 vccd1 _4192_/A sky130_fd_sc_hd__and4_2
XFILLER_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6558_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6845__105 vssd1 vssd1 vccd1 vccd1 _6845__105/HI _6954_/A sky130_fd_sc_hd__conb_1
XFILLER_105_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3520_ _6648_/Q _3534_/B _3516_/D _6649_/Q vssd1 vssd1 vccd1 vccd1 _3521_/D sky130_fd_sc_hd__a22o_1
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3451_ _6305_/Q _6509_/Q _3451_/S vssd1 vssd1 vccd1 vccd1 _3452_/A sky130_fd_sc_hd__mux2_1
X_3382_ _5412_/B _3385_/D _3382_/C vssd1 vssd1 vccd1 vccd1 _3383_/A sky130_fd_sc_hd__and3_1
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6170_ _6182_/B vssd1 vssd1 vccd1 vccd1 _6180_/B sky130_fd_sc_hd__clkbuf_1
X_5121_ _5119_/X _5120_/X _5115_/X vssd1 vssd1 vccd1 vccd1 _5122_/C sky130_fd_sc_hd__a21o_1
XFILLER_111_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _5086_/A vssd1 vssd1 vccd1 vccd1 _5181_/A sky130_fd_sc_hd__buf_2
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4003_ _4228_/A _4039_/C _4039_/D _4151_/A vssd1 vssd1 vccd1 vccd1 _4006_/A sky130_fd_sc_hd__a22oi_1
XFILLER_65_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5954_ _5935_/X _5952_/X _5953_/X _5687_/X vssd1 vssd1 vccd1 vccd1 _5954_/X sky130_fd_sc_hd__a211o_1
X_4905_ _4928_/A vssd1 vssd1 vccd1 vccd1 _4919_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5885_ _5935_/A _5885_/B vssd1 vssd1 vccd1 vccd1 _5885_/X sky130_fd_sc_hd__and2_1
XFILLER_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4836_ _4847_/A vssd1 vssd1 vccd1 vccd1 _4845_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_21_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4767_ _6402_/Q _4767_/B vssd1 vssd1 vccd1 vccd1 _4768_/A sky130_fd_sc_hd__and2_1
X_6506_ _6509_/CLK _6506_/D vssd1 vssd1 vccd1 vccd1 _6506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3718_ _3667_/X _3678_/Y _3708_/Y _3709_/X vssd1 vssd1 vccd1 vccd1 _3718_/X sky130_fd_sc_hd__a211o_1
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4698_ _6363_/Q _4700_/B vssd1 vssd1 vccd1 vccd1 _4699_/A sky130_fd_sc_hd__and2_1
XFILLER_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6437_ _6795_/CLK _6437_/D vssd1 vssd1 vccd1 vccd1 _6437_/Q sky130_fd_sc_hd__dfxtp_1
X_3649_ _3648_/B _3648_/C _3648_/A vssd1 vssd1 vccd1 vccd1 _3656_/C sky130_fd_sc_hd__a21o_1
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6368_ _6763_/CLK _6368_/D vssd1 vssd1 vccd1 vccd1 _6368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5319_ _5786_/C _5775_/B vssd1 vssd1 vccd1 vccd1 _5880_/B sky130_fd_sc_hd__nor2_1
XFILLER_102_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6299_ _6504_/CLK _6299_/D vssd1 vssd1 vccd1 vccd1 _6299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 _3330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5670_ _5670_/A _5670_/B vssd1 vssd1 vccd1 vccd1 _5670_/X sky130_fd_sc_hd__or2_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4621_ _4598_/A _4598_/B _4596_/B vssd1 vssd1 vccd1 vccd1 _4627_/A sky130_fd_sc_hd__o21ai_2
X_4552_ _4552_/A _4552_/B vssd1 vssd1 vccd1 vccd1 _4554_/A sky130_fd_sc_hd__xnor2_1
X_4483_ _4483_/A _4483_/B _4483_/C vssd1 vssd1 vccd1 vccd1 _4485_/B sky130_fd_sc_hd__nand3_1
X_3503_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3639_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6222_ _6286_/A _6222_/B vssd1 vssd1 vccd1 vccd1 _6222_/X sky130_fd_sc_hd__or2_1
X_3434_ _5214_/C _6505_/Q _3451_/S vssd1 vssd1 vccd1 vccd1 _3435_/A sky130_fd_sc_hd__mux2_1
X_3365_ _6551_/Q _6550_/Q _6332_/Q vssd1 vssd1 vccd1 vccd1 _4993_/C sky130_fd_sc_hd__nor3b_1
X_6153_ _6771_/Q _6142_/X _6151_/X _6152_/X vssd1 vssd1 vccd1 vccd1 _6771_/D sky130_fd_sc_hd__o211a_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5104_ _6813_/Q _5109_/B vssd1 vssd1 vccd1 vccd1 _5104_/X sky130_fd_sc_hd__or2_1
XFILLER_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3296_ _3298_/A vssd1 vssd1 vccd1 vccd1 _3296_/Y sky130_fd_sc_hd__inv_2
X_6084_ _6084_/A _6084_/B vssd1 vssd1 vccd1 vccd1 _6085_/A sky130_fd_sc_hd__and2_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5035_ _6895_/A _4945_/X _5033_/X _5034_/X vssd1 vssd1 vccd1 vccd1 _6557_/D sky130_fd_sc_hd__o211a_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6986_ _6986_/A _3291_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5937_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5957_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5868_ _5777_/X _5866_/X _5867_/Y _6493_/Q _5538_/X vssd1 vssd1 vccd1 vccd1 _5868_/X
+ sky130_fd_sc_hd__a221o_1
X_4819_ _6425_/Q _4823_/B vssd1 vssd1 vccd1 vccd1 _4820_/A sky130_fd_sc_hd__and2_1
X_5799_ _5542_/X _5798_/X _5814_/S vssd1 vssd1 vccd1 vccd1 _5799_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6771_ _6789_/CLK _6771_/D vssd1 vssd1 vccd1 vccd1 _6771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5722_ _6250_/A _5678_/X _5680_/X _5721_/X _5695_/X vssd1 vssd1 vccd1 vccd1 _5722_/X
+ sky130_fd_sc_hd__a221o_1
X_3983_ _3995_/A _3995_/B vssd1 vssd1 vccd1 vccd1 _4024_/B sky130_fd_sc_hd__xnor2_1
XFILLER_31_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5653_ _6685_/Q _5652_/X _5661_/S vssd1 vssd1 vccd1 vccd1 _5654_/B sky130_fd_sc_hd__mux2_1
X_4604_ _4605_/A _4605_/B vssd1 vssd1 vccd1 vccd1 _4606_/A sky130_fd_sc_hd__and2_1
X_5584_ _6452_/Q _5660_/B vssd1 vssd1 vccd1 vccd1 _5584_/X sky130_fd_sc_hd__and2_2
X_4535_ _4535_/A _4535_/B _4535_/C vssd1 vssd1 vccd1 vccd1 _4566_/D sky130_fd_sc_hd__and3_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4466_ _4466_/A vssd1 vssd1 vccd1 vccd1 _4466_/Y sky130_fd_sc_hd__inv_2
X_4397_ _6670_/Q vssd1 vssd1 vccd1 vccd1 _4576_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6205_ _6260_/A _6205_/B vssd1 vssd1 vccd1 vccd1 _6205_/X sky130_fd_sc_hd__or2_1
X_3417_ _3534_/B vssd1 vssd1 vccd1 vccd1 _5217_/B sky130_fd_sc_hd__clkbuf_2
X_3348_ _6328_/Q _3347_/Y _6330_/D vssd1 vssd1 vccd1 vccd1 _6328_/D sky130_fd_sc_hd__a21o_1
X_6136_ _6136_/A _6136_/B vssd1 vssd1 vccd1 vccd1 _6137_/A sky130_fd_sc_hd__and2_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _6067_/A _6067_/B vssd1 vssd1 vccd1 vccd1 _6752_/D sky130_fd_sc_hd__nor2_1
X_3279_ _3280_/A vssd1 vssd1 vccd1 vccd1 _3279_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5018_ _5176_/A vssd1 vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__buf_4
XFILLER_54_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6969_ _6969_/A _3271_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4320_ _4320_/A _4320_/B vssd1 vssd1 vccd1 vccd1 _4320_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4251_ _4249_/X _4238_/X _4240_/Y _4385_/A vssd1 vssd1 vccd1 vccd1 _4252_/B sky130_fd_sc_hd__a31o_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3202_ _3206_/A vssd1 vssd1 vccd1 vccd1 _3202_/Y sky130_fd_sc_hd__inv_2
X_4182_ _4202_/A _4058_/B _4183_/C vssd1 vssd1 vccd1 vccd1 _4184_/A sky130_fd_sc_hd__a21oi_1
XFILLER_95_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6754_ _6799_/CLK _6754_/D vssd1 vssd1 vccd1 vccd1 _6754_/Q sky130_fd_sc_hd__dfxtp_1
X_3966_ _4013_/A _4151_/B vssd1 vssd1 vccd1 vccd1 _3967_/B sky130_fd_sc_hd__nand2_1
X_6685_ _6532_/Q _6685_/D vssd1 vssd1 vccd1 vccd1 _6685_/Q sky130_fd_sc_hd__dfxtp_1
X_5705_ _5915_/A vssd1 vssd1 vccd1 vccd1 _5705_/X sky130_fd_sc_hd__clkbuf_2
X_5636_ _5630_/X _5631_/X _5620_/X _5635_/X vssd1 vssd1 vccd1 vccd1 _5636_/X sky130_fd_sc_hd__o211a_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3897_ _4103_/A _4257_/A _4262_/A _3889_/A vssd1 vssd1 vccd1 vccd1 _3899_/B sky130_fd_sc_hd__a22o_1
X_5567_ _6003_/A vssd1 vssd1 vccd1 vccd1 _5567_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4518_ _4518_/A _4518_/B vssd1 vssd1 vccd1 vccd1 _4541_/A sky130_fd_sc_hd__or2_1
X_5498_ _5498_/A vssd1 vssd1 vccd1 vccd1 _6671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4449_ _4449_/A _4545_/D vssd1 vssd1 vccd1 vccd1 _4453_/A sky130_fd_sc_hd__nand2_1
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6119_ _6762_/Q _6106_/X _6118_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6120_/B sky130_fd_sc_hd__a22o_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3820_ _3820_/A _3820_/B vssd1 vssd1 vccd1 vccd1 _3820_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3751_ _3751_/A _3751_/B vssd1 vssd1 vccd1 vccd1 _3751_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6470_ _6763_/CLK _6470_/D vssd1 vssd1 vccd1 vccd1 _6470_/Q sky130_fd_sc_hd__dfxtp_1
X_3682_ _6653_/Q _3720_/C vssd1 vssd1 vccd1 vccd1 _3684_/A sky130_fd_sc_hd__and2_1
X_5421_ _5217_/C _3706_/A _5431_/S vssd1 vssd1 vccd1 vccd1 _5422_/B sky130_fd_sc_hd__mux2_1
X_5352_ _5352_/A vssd1 vssd1 vccd1 vccd1 _6627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4303_ _4304_/B _4304_/C _4304_/A vssd1 vssd1 vccd1 vccd1 _4305_/B sky130_fd_sc_hd__o21ai_1
X_5283_ _5283_/A vssd1 vssd1 vccd1 vccd1 _6606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4234_ _4247_/B _4234_/B vssd1 vssd1 vccd1 vccd1 _4235_/B sky130_fd_sc_hd__xnor2_2
X_4165_ _4135_/B _4169_/B _4218_/A _4164_/X vssd1 vssd1 vccd1 vccd1 _4218_/B sky130_fd_sc_hd__a211oi_2
XFILLER_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4096_ _4135_/A _4096_/B vssd1 vssd1 vccd1 vccd1 _4098_/A sky130_fd_sc_hd__nor2_1
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6806_ _6809_/CLK _6806_/D vssd1 vssd1 vccd1 vccd1 _6806_/Q sky130_fd_sc_hd__dfxtp_1
X_4998_ _6549_/Q _4998_/B vssd1 vssd1 vccd1 vccd1 _4999_/C sky130_fd_sc_hd__nand2_1
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6737_ _6809_/CLK _6737_/D vssd1 vssd1 vccd1 vccd1 _6737_/Q sky130_fd_sc_hd__dfxtp_1
X_3949_ _3921_/Y _3936_/B _3927_/B _3927_/A vssd1 vssd1 vccd1 vccd1 _3951_/B sky130_fd_sc_hd__o22a_1
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6668_ _6795_/CLK _6668_/D vssd1 vssd1 vccd1 vccd1 _6668_/Q sky130_fd_sc_hd__dfxtp_1
X_6599_ _6667_/CLK _6599_/D vssd1 vssd1 vccd1 vccd1 _6599_/Q sky130_fd_sc_hd__dfxtp_1
X_5619_ _6472_/Q vssd1 vssd1 vccd1 vccd1 _5619_/X sky130_fd_sc_hd__buf_2
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5970_ _6635_/Q _6634_/Q _6633_/Q _6628_/Q vssd1 vssd1 vccd1 vccd1 _5972_/A sky130_fd_sc_hd__or4_2
XFILLER_52_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4921_ _4921_/A vssd1 vssd1 vccd1 vccd1 _6528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4852_ _6440_/Q _4856_/B vssd1 vssd1 vccd1 vccd1 _4853_/A sky130_fd_sc_hd__and2_1
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3803_ _3826_/A _3803_/B vssd1 vssd1 vccd1 vccd1 _3828_/D sky130_fd_sc_hd__xor2_2
X_4783_ _6409_/Q _4789_/B vssd1 vssd1 vccd1 vccd1 _4784_/A sky130_fd_sc_hd__and2_1
X_6522_ _6522_/CLK _6522_/D vssd1 vssd1 vccd1 vccd1 _6522_/Q sky130_fd_sc_hd__dfxtp_1
X_3734_ _3734_/A _3734_/B _3734_/C vssd1 vssd1 vccd1 vccd1 _3750_/B sky130_fd_sc_hd__nand3_2
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3665_ _3665_/A _3665_/B _3665_/C vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__and3_1
X_6453_ _6789_/CLK _6453_/D vssd1 vssd1 vccd1 vccd1 _6453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5404_ _3352_/X _5650_/A _5406_/B vssd1 vssd1 vccd1 vccd1 _5405_/B sky130_fd_sc_hd__mux2_1
X_6384_ _6795_/CLK _6384_/D vssd1 vssd1 vccd1 vccd1 _6384_/Q sky130_fd_sc_hd__dfxtp_1
X_3596_ _3596_/A _3722_/B _3596_/C vssd1 vssd1 vccd1 vccd1 _3596_/X sky130_fd_sc_hd__and3_1
XFILLER_88_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5335_ _6248_/A _5335_/B vssd1 vssd1 vccd1 vccd1 _5335_/X sky130_fd_sc_hd__or2_1
X_5266_ _5266_/A vssd1 vssd1 vccd1 vccd1 _6598_/D sky130_fd_sc_hd__clkbuf_1
X_4217_ _4239_/A _4217_/B vssd1 vssd1 vccd1 vccd1 _4217_/Y sky130_fd_sc_hd__nand2_1
X_5197_ _5243_/A _5197_/B _5197_/C vssd1 vssd1 vccd1 vccd1 _5198_/A sky130_fd_sc_hd__and3_1
XFILLER_56_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4148_ _4177_/A _4183_/B _4101_/A _4149_/B vssd1 vssd1 vccd1 vccd1 _4150_/A sky130_fd_sc_hd__a22oi_1
XFILLER_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4079_ _4079_/A _4079_/B _4079_/C vssd1 vssd1 vccd1 vccd1 _4081_/B sky130_fd_sc_hd__nand3_1
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6884__144 vssd1 vssd1 vccd1 vccd1 _6884__144/HI _6993_/A sky130_fd_sc_hd__conb_1
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3450_ _3450_/A vssd1 vssd1 vccd1 vccd1 _6304_/D sky130_fd_sc_hd__clkbuf_1
X_3381_ _6289_/Q _6290_/Q vssd1 vssd1 vccd1 vccd1 _3382_/C sky130_fd_sc_hd__or2_1
X_5120_ _6688_/Q _6720_/Q _6752_/Q _6784_/Q _4950_/B _4950_/A vssd1 vssd1 vccd1 vccd1
+ _5120_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5051_ _5077_/A _5051_/B vssd1 vssd1 vccd1 vccd1 _5051_/X sky130_fd_sc_hd__or2_1
XFILLER_111_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4002_ _4153_/B vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5953_ _6491_/Q _5957_/B _5957_/C vssd1 vssd1 vccd1 vccd1 _5953_/X sky130_fd_sc_hd__and3_1
XFILLER_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5884_ _6463_/Q _5919_/A _5890_/A _5941_/A _6721_/Q vssd1 vssd1 vccd1 vccd1 _5885_/B
+ sky130_fd_sc_hd__a32o_1
X_4904_ _6523_/Q _4870_/A _4873_/A input51/X vssd1 vssd1 vccd1 vccd1 _6523_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4835_ _4835_/A vssd1 vssd1 vccd1 vccd1 _6480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4766_ _4766_/A vssd1 vssd1 vccd1 vccd1 _6449_/D sky130_fd_sc_hd__clkbuf_1
X_3717_ _3717_/A vssd1 vssd1 vccd1 vccd1 _6342_/D sky130_fd_sc_hd__clkbuf_1
X_6505_ _6509_/CLK _6505_/D vssd1 vssd1 vccd1 vccd1 _6505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4697_ _4697_/A vssd1 vssd1 vccd1 vccd1 _6418_/D sky130_fd_sc_hd__clkbuf_1
X_6868__128 vssd1 vssd1 vccd1 vccd1 _6868__128/HI _6977_/A sky130_fd_sc_hd__conb_1
X_6436_ _6795_/CLK _6436_/D vssd1 vssd1 vccd1 vccd1 _6436_/Q sky130_fd_sc_hd__dfxtp_1
X_3648_ _3648_/A _3648_/B _3648_/C vssd1 vssd1 vccd1 vccd1 _3656_/B sky130_fd_sc_hd__nand3_1
X_3579_ _6651_/Q _6298_/Q _6297_/Q _6652_/Q vssd1 vssd1 vccd1 vccd1 _3585_/B sky130_fd_sc_hd__a22o_1
X_6367_ _6763_/CLK _6367_/D vssd1 vssd1 vccd1 vccd1 _6367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5318_ _6627_/Q _6626_/Q _6625_/Q vssd1 vssd1 vccd1 vccd1 _5775_/B sky130_fd_sc_hd__or3_4
XFILLER_102_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6298_ _6504_/CLK _6298_/D vssd1 vssd1 vccd1 vccd1 _6298_/Q sky130_fd_sc_hd__dfxtp_1
X_5249_ _6591_/Q _5249_/B vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__and2_1
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4609_/B _4620_/B vssd1 vssd1 vccd1 vccd1 _4630_/A sky130_fd_sc_hd__and2b_1
XFILLER_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4551_ _4551_/A _4551_/B vssd1 vssd1 vccd1 vccd1 _4552_/B sky130_fd_sc_hd__nor2_1
X_4482_ _4483_/B _4483_/C _4483_/A vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__a21o_1
X_3502_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3659_/A sky130_fd_sc_hd__clkbuf_2
X_6221_ _6798_/Q _6207_/A _6220_/X _6216_/X vssd1 vssd1 vccd1 vccd1 _6798_/D sky130_fd_sc_hd__o211a_1
X_3433_ _3499_/S vssd1 vssd1 vccd1 vccd1 _3451_/S sky130_fd_sc_hd__clkbuf_2
X_6152_ _6178_/A vssd1 vssd1 vccd1 vccd1 _6152_/X sky130_fd_sc_hd__buf_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3364_ _3361_/X _3363_/X _3340_/X vssd1 vssd1 vccd1 vccd1 _6333_/D sky130_fd_sc_hd__o21a_1
X_5103_ _5108_/A _5103_/B vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__or2_1
XFILLER_58_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3295_ _3298_/A vssd1 vssd1 vccd1 vccd1 _3295_/Y sky130_fd_sc_hd__inv_2
X_6083_ _6755_/Q _6080_/X _6082_/X _6076_/X vssd1 vssd1 vccd1 vccd1 _6084_/B sky130_fd_sc_hd__a22o_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _6136_/A vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__buf_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6985_ _6985_/A _3290_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
XFILLER_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5936_ _5619_/X _5919_/X _5920_/X _5912_/X _6730_/Q vssd1 vssd1 vccd1 vccd1 _5936_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5867_ _5870_/B _6143_/B vssd1 vssd1 vccd1 vccd1 _5867_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4818_ _4818_/A vssd1 vssd1 vccd1 vccd1 _6472_/D sky130_fd_sc_hd__clkbuf_1
X_5798_ _6706_/Q _5544_/X _5813_/S vssd1 vssd1 vccd1 vccd1 _5798_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4749_ _4749_/A vssd1 vssd1 vccd1 vccd1 _6441_/D sky130_fd_sc_hd__clkbuf_1
X_6419_ _6763_/CLK _6419_/D vssd1 vssd1 vccd1 vccd1 _6419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6770_ _6789_/CLK _6770_/D vssd1 vssd1 vccd1 vccd1 _6770_/Q sky130_fd_sc_hd__dfxtp_1
X_3982_ _4009_/A _3982_/B vssd1 vssd1 vccd1 vccd1 _3995_/B sky130_fd_sc_hd__nor2_1
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5721_ _5570_/X _5720_/X _5721_/S vssd1 vssd1 vccd1 vccd1 _5721_/X sky130_fd_sc_hd__mux2_1
X_5652_ _6459_/Q _5652_/B vssd1 vssd1 vccd1 vccd1 _5652_/X sky130_fd_sc_hd__and2_2
X_4603_ _4574_/A _4637_/B _4583_/B _4602_/X vssd1 vssd1 vccd1 vccd1 _4605_/B sky130_fd_sc_hd__a31oi_1
X_5583_ _5632_/A vssd1 vssd1 vccd1 vccd1 _5624_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4534_ _4535_/B _4535_/C _4535_/A vssd1 vssd1 vccd1 vccd1 _4566_/C sky130_fd_sc_hd__a21oi_2
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4465_ _4462_/X _4463_/Y _4464_/Y vssd1 vssd1 vccd1 vccd1 _6389_/D sky130_fd_sc_hd__o21a_1
X_4396_ _4519_/A _4512_/B _4396_/C _4450_/A vssd1 vssd1 vccd1 vccd1 _4450_/B sky130_fd_sc_hd__nand4_2
X_3416_ _3720_/D vssd1 vssd1 vccd1 vccd1 _3534_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6204_ _6791_/Q _6194_/X _6202_/X _6203_/X vssd1 vssd1 vccd1 vccd1 _6791_/D sky130_fd_sc_hd__o211a_1
X_3347_ _3347_/A _3347_/B vssd1 vssd1 vccd1 vccd1 _3347_/Y sky130_fd_sc_hd__nor2_1
X_6135_ _6766_/Q _6106_/A _6134_/X _5406_/C vssd1 vssd1 vccd1 vccd1 _6136_/B sky130_fd_sc_hd__a22o_1
XFILLER_58_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6066_ _6752_/Q _6061_/X _6065_/X vssd1 vssd1 vccd1 vccd1 _6067_/B sky130_fd_sc_hd__a21oi_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _3280_/A vssd1 vssd1 vccd1 vccd1 _3278_/Y sky130_fd_sc_hd__inv_2
X_5017_ _5017_/A _5017_/B _5017_/C vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__nand3_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6968_ _6968_/A _3270_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5919_ _5919_/A vssd1 vssd1 vccd1 vccd1 _5919_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6899_ _6899_/A _3186_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__ebufn_8
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4250_ _4238_/X _4240_/Y _4249_/X vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__a21oi_1
XFILLER_4_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3201_ _3219_/A vssd1 vssd1 vccd1 vccd1 _3206_/A sky130_fd_sc_hd__buf_2
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4181_ _4181_/A _4205_/A vssd1 vssd1 vccd1 vccd1 _4183_/C sky130_fd_sc_hd__nor2_1
XFILLER_79_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6753_ _6799_/CLK _6753_/D vssd1 vssd1 vccd1 vccd1 _6753_/Q sky130_fd_sc_hd__dfxtp_1
X_3965_ _4180_/D vssd1 vssd1 vccd1 vccd1 _4151_/B sky130_fd_sc_hd__buf_2
X_6684_ _6532_/Q _6684_/D vssd1 vssd1 vccd1 vccd1 _6684_/Q sky130_fd_sc_hd__dfxtp_1
X_5704_ _5734_/A vssd1 vssd1 vccd1 vccd1 _5704_/X sky130_fd_sc_hd__clkbuf_2
X_3896_ _4039_/D vssd1 vssd1 vccd1 vccd1 _4262_/A sky130_fd_sc_hd__clkbuf_2
X_5635_ _5670_/A _5635_/B vssd1 vssd1 vccd1 vccd1 _5635_/X sky130_fd_sc_hd__or2_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5566_ _6031_/A vssd1 vssd1 vccd1 vccd1 _6003_/A sky130_fd_sc_hd__buf_2
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4517_ _4517_/A _4517_/B _6379_/Q _6380_/Q vssd1 vssd1 vccd1 vccd1 _4518_/B sky130_fd_sc_hd__and4_1
X_5497_ _6084_/A _5497_/B vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__and2_1
X_4448_ _6381_/Q vssd1 vssd1 vccd1 vccd1 _4545_/D sky130_fd_sc_hd__buf_2
XFILLER_120_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _4379_/A _4379_/B vssd1 vssd1 vccd1 vccd1 _4381_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6118_ _6472_/Q _6107_/X _6096_/X _6113_/X _6488_/Q vssd1 vssd1 vccd1 vccd1 _6118_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6492_/Q _6023_/A _6249_/A _6031_/X vssd1 vssd1 vccd1 vccd1 _6049_/X sky130_fd_sc_hd__a31o_1
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3750_ _3750_/A _3750_/B _3750_/C vssd1 vssd1 vccd1 vccd1 _3750_/Y sky130_fd_sc_hd__nand3_1
XFILLER_20_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3681_ _3789_/A _3789_/B _3720_/D _3681_/D vssd1 vssd1 vccd1 vccd1 _3684_/C sky130_fd_sc_hd__nand4_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5420_ _5420_/A vssd1 vssd1 vccd1 vccd1 _6648_/D sky130_fd_sc_hd__clkbuf_1
X_5351_ _6627_/Q _5372_/B vssd1 vssd1 vccd1 vccd1 _5352_/A sky130_fd_sc_hd__and2_1
XFILLER_114_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5282_ _6606_/Q _5282_/B vssd1 vssd1 vccd1 vccd1 _5283_/A sky130_fd_sc_hd__and2_1
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4302_ _4333_/A _4300_/B _4301_/Y _4296_/X vssd1 vssd1 vccd1 vccd1 _4304_/C sky130_fd_sc_hd__o2bb2a_1
XFILLER_102_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4233_ _4243_/A _4247_/A vssd1 vssd1 vccd1 vccd1 _4234_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4164_ _4176_/B _4162_/Y _4144_/B _4144_/Y vssd1 vssd1 vccd1 vccd1 _4164_/X sky130_fd_sc_hd__o211a_1
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4095_ _3992_/A _4101_/A _4049_/B _4093_/Y vssd1 vssd1 vccd1 vccd1 _4096_/B sky130_fd_sc_hd__a211oi_1
XFILLER_83_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6805_ _6809_/CLK _6805_/D vssd1 vssd1 vccd1 vccd1 _6805_/Q sky130_fd_sc_hd__dfxtp_1
X_4997_ _6549_/Q _4998_/B vssd1 vssd1 vccd1 vccd1 _4999_/B sky130_fd_sc_hd__or2_1
X_6736_ _6809_/CLK _6736_/D vssd1 vssd1 vccd1 vccd1 _6736_/Q sky130_fd_sc_hd__dfxtp_1
X_3948_ _3959_/A _3959_/B vssd1 vssd1 vccd1 vccd1 _3951_/A sky130_fd_sc_hd__xnor2_1
X_6667_ _6667_/CLK _6667_/D vssd1 vssd1 vccd1 vccd1 _6667_/Q sky130_fd_sc_hd__dfxtp_1
X_3879_ _3879_/A _4257_/B vssd1 vssd1 vccd1 vccd1 _3880_/A sky130_fd_sc_hd__and2_1
X_6598_ _6667_/CLK _6598_/D vssd1 vssd1 vccd1 vccd1 _6598_/Q sky130_fd_sc_hd__dfxtp_1
X_5618_ _6681_/Q _5601_/X _5614_/X _5617_/X _5591_/X vssd1 vssd1 vccd1 vccd1 _6681_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5549_ _6237_/A _5534_/X _6286_/B _5538_/X vssd1 vssd1 vccd1 vccd1 _5549_/X sky130_fd_sc_hd__a31o_1
XFILLER_105_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6816__76 vssd1 vssd1 vccd1 vccd1 _6816__76/HI _6925_/A sky130_fd_sc_hd__conb_1
XFILLER_86_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ _4919_/X _6528_/Q _4926_/S vssd1 vssd1 vccd1 vccd1 _4921_/A sky130_fd_sc_hd__mux2_1
X_6830__90 vssd1 vssd1 vccd1 vccd1 _6830__90/HI _6939_/A sky130_fd_sc_hd__conb_1
X_4851_ _4851_/A vssd1 vssd1 vccd1 vccd1 _6487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3802_ _3806_/A _3806_/B vssd1 vssd1 vccd1 vccd1 _3803_/B sky130_fd_sc_hd__xnor2_2
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4782_ _4782_/A vssd1 vssd1 vccd1 vccd1 _6456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6521_ _6523_/CLK _6521_/D vssd1 vssd1 vccd1 vccd1 _6521_/Q sky130_fd_sc_hd__dfxtp_1
X_3733_ _3694_/A _3694_/C _3694_/B vssd1 vssd1 vccd1 vccd1 _3734_/C sky130_fd_sc_hd__a21bo_1
X_3664_ _3665_/B _3665_/C _3665_/A vssd1 vssd1 vccd1 vccd1 _3664_/Y sky130_fd_sc_hd__a21oi_1
X_6452_ _6789_/CLK _6452_/D vssd1 vssd1 vccd1 vccd1 _6452_/Q sky130_fd_sc_hd__dfxtp_1
X_5403_ _5403_/A vssd1 vssd1 vccd1 vccd1 _6643_/D sky130_fd_sc_hd__clkbuf_1
X_6383_ _6795_/CLK _6383_/D vssd1 vssd1 vccd1 vccd1 _6383_/Q sky130_fd_sc_hd__dfxtp_1
X_3595_ _3595_/A vssd1 vssd1 vccd1 vccd1 _6339_/D sky130_fd_sc_hd__clkbuf_1
X_5334_ _6268_/A vssd1 vssd1 vccd1 vccd1 _6248_/A sky130_fd_sc_hd__clkbuf_4
X_5265_ _6598_/Q _5271_/B vssd1 vssd1 vccd1 vccd1 _5266_/A sky130_fd_sc_hd__and2_1
XFILLER_102_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5196_ _5181_/X _5195_/X _5176_/X vssd1 vssd1 vccd1 vccd1 _5197_/C sky130_fd_sc_hd__a21o_1
X_4216_ _4216_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _4217_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4147_ _4147_/A vssd1 vssd1 vccd1 vccd1 _4177_/A sky130_fd_sc_hd__buf_2
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4078_ _4079_/B _4079_/C _4079_/A vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__a21o_1
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6719_ _6809_/CLK _6719_/D vssd1 vssd1 vccd1 vccd1 _6719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3380_ _6289_/Q _6290_/Q vssd1 vssd1 vccd1 vccd1 _3385_/D sky130_fd_sc_hd__nand2_1
XFILLER_123_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5050_ _6677_/Q _6709_/Q _6741_/Q _6773_/Q _5049_/X _5029_/X vssd1 vssd1 vccd1 vccd1
+ _5051_/B sky130_fd_sc_hd__mux4_1
XFILLER_111_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4001_ _6662_/Q vssd1 vssd1 vccd1 vccd1 _4153_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5952_ _5651_/X _5947_/X _5920_/A _5961_/B _6733_/Q vssd1 vssd1 vccd1 vccd1 _5952_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4903_ _6522_/Q _4870_/A _4873_/A input50/X vssd1 vssd1 vccd1 vccd1 _6522_/D sky130_fd_sc_hd__a22o_1
X_5883_ _6107_/A vssd1 vssd1 vccd1 vccd1 _5919_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4834_ _6432_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4835_/A sky130_fd_sc_hd__and2_1
X_4765_ _6401_/Q _4767_/B vssd1 vssd1 vccd1 vccd1 _4766_/A sky130_fd_sc_hd__and2_1
XFILLER_119_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3716_ _3899_/A _3716_/B _3716_/C vssd1 vssd1 vccd1 vccd1 _3717_/A sky130_fd_sc_hd__and3_1
X_6504_ _6504_/CLK _6504_/D vssd1 vssd1 vccd1 vccd1 _6504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4696_ _6362_/Q _4700_/B vssd1 vssd1 vccd1 vccd1 _4697_/A sky130_fd_sc_hd__and2_1
X_6435_ _6795_/CLK _6435_/D vssd1 vssd1 vccd1 vccd1 _6435_/Q sky130_fd_sc_hd__dfxtp_1
X_3647_ _3647_/A _3647_/B _3647_/C vssd1 vssd1 vccd1 vccd1 _3648_/C sky130_fd_sc_hd__nand3_1
X_3578_ _3757_/A _3578_/B vssd1 vssd1 vccd1 vccd1 _3586_/A sky130_fd_sc_hd__nand2_1
X_6366_ _6763_/CLK _6366_/D vssd1 vssd1 vccd1 vccd1 _6366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5317_ _6620_/Q vssd1 vssd1 vccd1 vccd1 _5786_/C sky130_fd_sc_hd__inv_2
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6297_ _6504_/CLK _6297_/D vssd1 vssd1 vccd1 vccd1 _6297_/Q sky130_fd_sc_hd__dfxtp_1
X_5248_ _5248_/A vssd1 vssd1 vccd1 vccd1 _6590_/D sky130_fd_sc_hd__clkbuf_1
X_5179_ _5179_/A vssd1 vssd1 vccd1 vccd1 _6580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6851__111 vssd1 vssd1 vccd1 vccd1 _6851__111/HI _6960_/A sky130_fd_sc_hd__conb_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4550_ _4576_/A _4576_/B _4550_/C _4576_/C vssd1 vssd1 vccd1 vccd1 _4551_/B sky130_fd_sc_hd__and4_1
X_4481_ _4481_/A _4481_/B vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__xnor2_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3501_ _6648_/Q vssd1 vssd1 vccd1 vccd1 _3616_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6220_ _6283_/A _6222_/B vssd1 vssd1 vccd1 vccd1 _6220_/X sky130_fd_sc_hd__or2_1
X_3432_ _3808_/D vssd1 vssd1 vccd1 vccd1 _5214_/C sky130_fd_sc_hd__buf_2
X_3363_ _4980_/B _3362_/Y _6333_/Q vssd1 vssd1 vccd1 vccd1 _3363_/X sky130_fd_sc_hd__o21a_1
X_6151_ _6240_/A _6154_/B vssd1 vssd1 vccd1 vccd1 _6151_/X sky130_fd_sc_hd__or2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5102_ _6685_/Q _6717_/Q _6749_/Q _6781_/Q _5083_/X _4949_/A vssd1 vssd1 vccd1 vccd1
+ _5103_/B sky130_fd_sc_hd__mux4_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3294_ _3298_/A vssd1 vssd1 vccd1 vccd1 _3294_/Y sky130_fd_sc_hd__inv_2
X_6082_ _6465_/Q _6081_/X _6070_/X _6138_/S _6481_/Q vssd1 vssd1 vccd1 vccd1 _6082_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5033_ _5011_/X _5031_/X _5032_/X _5019_/X vssd1 vssd1 vccd1 vccd1 _5033_/X sky130_fd_sc_hd__a31o_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6984_ _6984_/A _3289_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5935_ _5935_/A vssd1 vssd1 vccd1 vccd1 _5935_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5866_ _6477_/Q _5865_/X _5866_/S vssd1 vssd1 vccd1 vccd1 _5866_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4817_ _6424_/Q _4823_/B vssd1 vssd1 vccd1 vccd1 _4818_/A sky130_fd_sc_hd__and2_1
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5797_ _5797_/A vssd1 vssd1 vccd1 vccd1 _5797_/X sky130_fd_sc_hd__clkbuf_2
X_4748_ _6393_/Q _4756_/B vssd1 vssd1 vccd1 vccd1 _4749_/A sky130_fd_sc_hd__and2_1
XFILLER_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4679_ _4679_/A vssd1 vssd1 vccd1 vccd1 _4688_/B sky130_fd_sc_hd__clkbuf_2
X_6418_ _6763_/CLK _6418_/D vssd1 vssd1 vccd1 vccd1 _6418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6349_ _6789_/CLK _6349_/D vssd1 vssd1 vccd1 vccd1 _6349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3981_ _4202_/A _3979_/D _3973_/X _3977_/X vssd1 vssd1 vccd1 vccd1 _3982_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5720_ _6693_/Q _5572_/X _5751_/S vssd1 vssd1 vccd1 vccd1 _5720_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5651_ _6475_/Q vssd1 vssd1 vccd1 vccd1 _5651_/X sky130_fd_sc_hd__buf_2
X_4602_ _4582_/B _4602_/B vssd1 vssd1 vccd1 vccd1 _4602_/X sky130_fd_sc_hd__and2b_1
X_5582_ _5631_/A vssd1 vssd1 vccd1 vccd1 _5582_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4533_ _4502_/A _4502_/C _4502_/B vssd1 vssd1 vccd1 vccd1 _4535_/A sky130_fd_sc_hd__a21bo_1
XFILLER_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4464_ _4462_/X _4463_/Y _3637_/A vssd1 vssd1 vccd1 vccd1 _4464_/Y sky130_fd_sc_hd__a21oi_1
X_6203_ _6255_/A vssd1 vssd1 vccd1 vccd1 _6203_/X sky130_fd_sc_hd__buf_2
X_4395_ _6378_/Q vssd1 vssd1 vccd1 vccd1 _4512_/B sky130_fd_sc_hd__buf_2
X_3415_ _6298_/Q vssd1 vssd1 vccd1 vccd1 _3720_/D sky130_fd_sc_hd__clkbuf_2
X_6134_ _6476_/Q _5919_/A _6070_/A _6113_/A _6492_/Q vssd1 vssd1 vccd1 vccd1 _6134_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_58_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3346_ _3346_/A _3346_/B _3346_/C vssd1 vssd1 vccd1 vccd1 _3347_/B sky130_fd_sc_hd__or3_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6065_ _6478_/Q _6058_/Y _6064_/X _5824_/A vssd1 vssd1 vccd1 vccd1 _6065_/X sky130_fd_sc_hd__o211a_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3277_ _3280_/A vssd1 vssd1 vccd1 vccd1 _3277_/Y sky130_fd_sc_hd__inv_2
X_5016_ _5015_/X _6800_/Q _5113_/A vssd1 vssd1 vccd1 vccd1 _5016_/X sky130_fd_sc_hd__mux2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6967_ _6967_/A _3268_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
X_5918_ _5946_/A vssd1 vssd1 vccd1 vccd1 _5918_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6898_ _6898_/A _3185_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__ebufn_8
X_5849_ _6715_/Q _5825_/X _5848_/X _5838_/X vssd1 vssd1 vccd1 vccd1 _6715_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3200_ _3200_/A vssd1 vssd1 vccd1 vccd1 _3200_/Y sky130_fd_sc_hd__inv_2
X_4180_ _4227_/A _4180_/B _4180_/C _4180_/D vssd1 vssd1 vccd1 vccd1 _4205_/A sky130_fd_sc_hd__and4_1
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6752_ _6799_/CLK _6752_/D vssd1 vssd1 vccd1 vccd1 _6752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3964_ _6355_/Q vssd1 vssd1 vccd1 vccd1 _4180_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6683_ _6532_/Q _6683_/D vssd1 vssd1 vccd1 vccd1 _6683_/Q sky130_fd_sc_hd__dfxtp_1
X_3895_ _4076_/C vssd1 vssd1 vccd1 vccd1 _4039_/D sky130_fd_sc_hd__clkbuf_2
X_5703_ _5542_/X _5698_/X _5699_/X _5702_/X vssd1 vssd1 vccd1 vccd1 _5703_/X sky130_fd_sc_hd__o211a_1
X_5634_ _6683_/Q _5633_/X _5661_/S vssd1 vssd1 vccd1 vccd1 _5635_/B sky130_fd_sc_hd__mux2_1
X_5565_ _6482_/Q vssd1 vssd1 vccd1 vccd1 _6243_/A sky130_fd_sc_hd__buf_2
X_4516_ _4517_/A _6379_/Q _6380_/Q _4517_/B vssd1 vssd1 vccd1 vccd1 _4518_/A sky130_fd_sc_hd__a22oi_1
X_5496_ _6319_/Q _4637_/A _5496_/S vssd1 vssd1 vccd1 vccd1 _5497_/B sky130_fd_sc_hd__mux2_1
X_4447_ _4468_/B _4468_/C _4468_/A vssd1 vssd1 vccd1 vccd1 _4455_/C sky130_fd_sc_hd__a21o_1
XFILLER_120_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4378_ _4418_/A _4418_/B vssd1 vssd1 vccd1 vccd1 _4379_/B sky130_fd_sc_hd__xor2_1
XFILLER_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6117_ _6117_/A vssd1 vssd1 vccd1 vccd1 _6761_/D sky130_fd_sc_hd__clkbuf_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3329_ _3329_/A _3329_/B _3329_/C _3329_/D vssd1 vssd1 vccd1 vccd1 _3329_/X sky130_fd_sc_hd__or4_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6048_ _6750_/Q _5659_/X _6048_/S vssd1 vssd1 vccd1 vccd1 _6048_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6569_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3680_ _3759_/A _3645_/B _3681_/D _6655_/Q vssd1 vssd1 vccd1 vccd1 _3684_/B sky130_fd_sc_hd__a22o_1
X_5350_ _5350_/A vssd1 vssd1 vccd1 vccd1 _6626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5281_ _5281_/A vssd1 vssd1 vccd1 vccd1 _6605_/D sky130_fd_sc_hd__clkbuf_1
X_4301_ _4301_/A vssd1 vssd1 vccd1 vccd1 _4301_/Y sky130_fd_sc_hd__clkinv_2
X_4232_ _4232_/A _4232_/B vssd1 vssd1 vccd1 vccd1 _4247_/B sky130_fd_sc_hd__xnor2_2
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4163_ _4144_/B _4144_/Y _4176_/B _4162_/Y vssd1 vssd1 vccd1 vccd1 _4218_/A sky130_fd_sc_hd__a211oi_4
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4094_ _4049_/B _4093_/Y _3992_/A _4101_/A vssd1 vssd1 vccd1 vccd1 _4135_/A sky130_fd_sc_hd__o211a_1
XFILLER_83_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4996_ _6548_/Q _4996_/B vssd1 vssd1 vccd1 vccd1 _4998_/B sky130_fd_sc_hd__and2_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6804_ _6809_/CLK _6804_/D vssd1 vssd1 vccd1 vccd1 _6804_/Q sky130_fd_sc_hd__dfxtp_1
X_6735_ _6809_/CLK _6735_/D vssd1 vssd1 vccd1 vccd1 _6735_/Q sky130_fd_sc_hd__dfxtp_1
X_3947_ _3947_/A _3947_/B vssd1 vssd1 vccd1 vccd1 _3959_/B sky130_fd_sc_hd__xnor2_2
XFILLER_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6666_ _6667_/CLK _6666_/D vssd1 vssd1 vccd1 vccd1 _6666_/Q sky130_fd_sc_hd__dfxtp_1
X_3878_ _3878_/A vssd1 vssd1 vccd1 vccd1 _6355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6597_ _6667_/CLK _6597_/D vssd1 vssd1 vccd1 vccd1 _6597_/Q sky130_fd_sc_hd__dfxtp_1
X_5617_ _6263_/A _5589_/X _5578_/X _5616_/X vssd1 vssd1 vccd1 vccd1 _5617_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5548_ _6480_/Q vssd1 vssd1 vccd1 vccd1 _6237_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5479_ _5479_/A vssd1 vssd1 vccd1 vccd1 _6665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4850_ _6439_/Q _4856_/B vssd1 vssd1 vccd1 vccd1 _4851_/A sky130_fd_sc_hd__and2_1
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3801_ _3801_/A _3801_/B vssd1 vssd1 vccd1 vccd1 _3806_/B sky130_fd_sc_hd__xnor2_2
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6520_ _6523_/CLK _6520_/D vssd1 vssd1 vccd1 vccd1 _6520_/Q sky130_fd_sc_hd__dfxtp_1
X_4781_ _6408_/Q _4789_/B vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__and2_1
X_3732_ _3769_/A _3752_/B _3730_/X vssd1 vssd1 vccd1 vccd1 _3734_/B sky130_fd_sc_hd__or3b_1
X_3663_ _3663_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3665_/A sky130_fd_sc_hd__xnor2_1
X_6451_ _6789_/CLK _6451_/D vssd1 vssd1 vccd1 vccd1 _6451_/Q sky130_fd_sc_hd__dfxtp_1
X_5402_ _6643_/Q _5412_/B vssd1 vssd1 vccd1 vccd1 _5403_/A sky130_fd_sc_hd__and2_1
X_6382_ _6795_/CLK _6382_/D vssd1 vssd1 vccd1 vccd1 _6382_/Q sky130_fd_sc_hd__dfxtp_1
X_5333_ _6622_/Q vssd1 vssd1 vccd1 vccd1 _6268_/A sky130_fd_sc_hd__clkbuf_2
X_3594_ _3592_/X _5008_/B _3594_/C vssd1 vssd1 vccd1 vccd1 _3595_/A sky130_fd_sc_hd__and3b_1
X_5264_ _5264_/A vssd1 vssd1 vccd1 vccd1 _6597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5195_ _6700_/Q _6732_/Q _6764_/Q _6796_/Q _5188_/X _5169_/X vssd1 vssd1 vccd1 vccd1
+ _5195_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4215_ _4216_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__or2_1
X_4146_ _4160_/A _4146_/B _4124_/X vssd1 vssd1 vccd1 vccd1 _4160_/B sky130_fd_sc_hd__nor3b_1
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _6661_/Q _6353_/Q vssd1 vssd1 vccd1 vccd1 _4079_/A sky130_fd_sc_hd__and2_1
XFILLER_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4979_ _3329_/X _4979_/B _4979_/C _4979_/D vssd1 vssd1 vccd1 vccd1 _5008_/C sky130_fd_sc_hd__and4b_1
X_6718_ _6799_/CLK _6718_/D vssd1 vssd1 vccd1 vccd1 _6718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6649_ _6763_/CLK _6649_/D vssd1 vssd1 vccd1 vccd1 _6649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4000_ _4083_/A _4116_/B _4000_/C _4057_/A vssd1 vssd1 vccd1 vccd1 _4057_/B sky130_fd_sc_hd__nand4_2
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5951_ _6732_/Q _5946_/X _5950_/X _5933_/X vssd1 vssd1 vccd1 vccd1 _6732_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4902_ _6521_/Q _4870_/A _4873_/A input49/X vssd1 vssd1 vccd1 vccd1 _6521_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5882_ _5882_/A _5882_/B vssd1 vssd1 vccd1 vccd1 _6107_/A sky130_fd_sc_hd__and2_2
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4833_ _4833_/A vssd1 vssd1 vccd1 vccd1 _6479_/D sky130_fd_sc_hd__clkbuf_1
X_4764_ _4764_/A vssd1 vssd1 vccd1 vccd1 _6448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3715_ _3715_/A _3828_/A vssd1 vssd1 vccd1 vccd1 _3716_/C sky130_fd_sc_hd__or2_1
X_6503_ _6504_/CLK _6503_/D vssd1 vssd1 vccd1 vccd1 _6503_/Q sky130_fd_sc_hd__dfxtp_1
X_6434_ _6795_/CLK _6434_/D vssd1 vssd1 vccd1 vccd1 _6434_/Q sky130_fd_sc_hd__dfxtp_1
X_4695_ _4695_/A vssd1 vssd1 vccd1 vccd1 _6417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3646_ _3647_/B _3647_/C _3647_/A vssd1 vssd1 vccd1 vccd1 _3648_/B sky130_fd_sc_hd__a21o_1
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3577_ _6653_/Q vssd1 vssd1 vccd1 vccd1 _3757_/A sky130_fd_sc_hd__clkbuf_2
X_6365_ _6763_/CLK _6365_/D vssd1 vssd1 vccd1 vccd1 _6365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5316_ _6623_/Q vssd1 vssd1 vccd1 vccd1 _6224_/A sky130_fd_sc_hd__clkbuf_2
X_6296_ _6504_/CLK _6296_/D vssd1 vssd1 vccd1 vccd1 _6296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5247_ _6590_/Q _5249_/B vssd1 vssd1 vccd1 vccd1 _5248_/A sky130_fd_sc_hd__and2_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5178_ _5191_/A _5178_/B _5178_/C vssd1 vssd1 vccd1 vccd1 _5179_/A sky130_fd_sc_hd__and3_1
XFILLER_56_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4129_ _4128_/A _4128_/B _4128_/C vssd1 vssd1 vccd1 vccd1 _4144_/C sky130_fd_sc_hd__a21o_1
XFILLER_44_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6890__150 vssd1 vssd1 vccd1 vccd1 _6890__150/HI _6999_/A sky130_fd_sc_hd__conb_1
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3500_ _3500_/A vssd1 vssd1 vccd1 vccd1 _6327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4480_ _4480_/A _4480_/B vssd1 vssd1 vccd1 vccd1 _4481_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3431_ _3758_/B vssd1 vssd1 vccd1 vccd1 _3808_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3362_ _4993_/A _5017_/A vssd1 vssd1 vccd1 vccd1 _3362_/Y sky130_fd_sc_hd__nand2_1
X_6150_ _6770_/Q _6142_/X _6149_/X _6051_/X vssd1 vssd1 vccd1 vccd1 _6770_/D sky130_fd_sc_hd__o211a_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _6905_/A _5075_/X _5099_/X _5100_/X vssd1 vssd1 vccd1 vccd1 _6567_/D sky130_fd_sc_hd__o211a_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3305_/A vssd1 vssd1 vccd1 vccd1 _3298_/A sky130_fd_sc_hd__buf_12
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6562_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_6081_ _6107_/A vssd1 vssd1 vccd1 vccd1 _6081_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5032_ _6802_/Q _5044_/B vssd1 vssd1 vccd1 vccd1 _5032_/X sky130_fd_sc_hd__or2_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6983_ _6983_/A _3288_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
X_5934_ _6729_/Q _5918_/X _5932_/X _5933_/X vssd1 vssd1 vccd1 vccd1 _6729_/D sky130_fd_sc_hd__o211a_1
X_6874__134 vssd1 vssd1 vccd1 vccd1 _6874__134/HI _6983_/A sky130_fd_sc_hd__conb_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5865_ _6719_/Q _5668_/X _5865_/S vssd1 vssd1 vccd1 vccd1 _5865_/X sky130_fd_sc_hd__mux2_1
X_4816_ _4816_/A vssd1 vssd1 vccd1 vccd1 _6471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5796_ _6705_/Q _5755_/X _5795_/X _5773_/X vssd1 vssd1 vccd1 vccd1 _6705_/D sky130_fd_sc_hd__o211a_1
X_4747_ _4791_/A vssd1 vssd1 vccd1 vccd1 _4756_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4678_ _4678_/A vssd1 vssd1 vccd1 vccd1 _6410_/D sky130_fd_sc_hd__clkbuf_1
X_3629_ _3629_/A _3629_/B _3629_/C vssd1 vssd1 vccd1 vccd1 _3629_/X sky130_fd_sc_hd__and3_1
X_6417_ _6763_/CLK _6417_/D vssd1 vssd1 vccd1 vccd1 _6417_/Q sky130_fd_sc_hd__dfxtp_1
X_6348_ _6789_/CLK _6348_/D vssd1 vssd1 vccd1 vccd1 _6348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6279_ _6812_/Q _6267_/X _6278_/Y _6275_/X vssd1 vssd1 vccd1 vccd1 _6812_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6858__118 vssd1 vssd1 vccd1 vccd1 _6858__118/HI _6967_/A sky130_fd_sc_hd__conb_1
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _4151_/A vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5650_ _5650_/A vssd1 vssd1 vccd1 vccd1 _5650_/X sky130_fd_sc_hd__buf_2
XFILLER_31_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4601_ _4638_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__or2_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5581_ _6468_/Q vssd1 vssd1 vccd1 vccd1 _5581_/X sky130_fd_sc_hd__clkbuf_4
X_4532_ _4531_/B _4531_/C _4531_/A vssd1 vssd1 vccd1 vccd1 _4535_/C sky130_fd_sc_hd__a21o_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4463_ _4463_/A _4463_/B vssd1 vssd1 vccd1 vccd1 _4463_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3414_ _3414_/A vssd1 vssd1 vccd1 vccd1 _6297_/D sky130_fd_sc_hd__clkbuf_1
X_6202_ _6257_/A _6205_/B vssd1 vssd1 vccd1 vccd1 _6202_/X sky130_fd_sc_hd__or2_1
XFILLER_98_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4394_ _4477_/A _4388_/B _4396_/C _4450_/A vssd1 vssd1 vccd1 vccd1 _4429_/A sky130_fd_sc_hd__a22o_1
X_6133_ _6133_/A vssd1 vssd1 vccd1 vccd1 _6765_/D sky130_fd_sc_hd__clkbuf_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _6449_/Q _6448_/Q _6447_/Q _6446_/Q vssd1 vssd1 vccd1 vccd1 _3346_/C sky130_fd_sc_hd__or4_1
X_3276_ _3280_/A vssd1 vssd1 vccd1 vccd1 _3276_/Y sky130_fd_sc_hd__inv_2
X_6064_ _5971_/A _5873_/A _6462_/Q _5971_/B _6138_/S vssd1 vssd1 vccd1 vccd1 _6064_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5015_ _6672_/Q _6704_/Q _6736_/Q _6768_/Q _5012_/X _5014_/X vssd1 vssd1 vccd1 vccd1
+ _5015_/X sky130_fd_sc_hd__mux4_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6966_ _6966_/A _3267_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5917_ _6726_/Q _5888_/X _5916_/X _5904_/X vssd1 vssd1 vccd1 vccd1 _6726_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6897_ _6897_/A _3184_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__ebufn_8
X_5848_ _6489_/Q _5840_/X _5847_/X _5836_/X _5843_/X vssd1 vssd1 vccd1 vccd1 _5848_/X
+ sky130_fd_sc_hd__a221o_1
X_5779_ _5865_/S vssd1 vssd1 vccd1 vccd1 _5859_/S sky130_fd_sc_hd__buf_2
XFILLER_89_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6837__97 vssd1 vssd1 vccd1 vccd1 _6837__97/HI _6946_/A sky130_fd_sc_hd__conb_1
XFILLER_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6751_ _6799_/CLK _6751_/D vssd1 vssd1 vccd1 vccd1 _6751_/Q sky130_fd_sc_hd__dfxtp_1
X_3963_ _3992_/C _3963_/B vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_6682_ _6532_/Q _6682_/D vssd1 vssd1 vccd1 vccd1 _6682_/Q sky130_fd_sc_hd__dfxtp_1
X_3894_ _6351_/Q vssd1 vssd1 vccd1 vccd1 _4076_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5702_ _5765_/A _5702_/B vssd1 vssd1 vccd1 vccd1 _5702_/X sky130_fd_sc_hd__or2_1
X_5633_ _6457_/Q _5652_/B vssd1 vssd1 vccd1 vccd1 _5633_/X sky130_fd_sc_hd__and2_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5564_ _5560_/X _5525_/X _5505_/X _5563_/X vssd1 vssd1 vccd1 vccd1 _5564_/X sky130_fd_sc_hd__o211a_1
X_4515_ _4514_/A _4553_/B _4514_/C vssd1 vssd1 vccd1 vccd1 _4542_/B sky130_fd_sc_hd__a21oi_1
XFILLER_105_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5495_ _5495_/A vssd1 vssd1 vccd1 vccd1 _6670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4446_ _4468_/A _4468_/B _4468_/C vssd1 vssd1 vccd1 vccd1 _4455_/B sky130_fd_sc_hd__nand3_1
X_4377_ _4390_/A _4390_/B vssd1 vssd1 vccd1 vccd1 _4418_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6116_ _6132_/A _6116_/B vssd1 vssd1 vccd1 vccd1 _6117_/A sky130_fd_sc_hd__and2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ input7/X input6/X input9/X input8/X vssd1 vssd1 vccd1 vccd1 _3329_/D sky130_fd_sc_hd__or4_2
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _3262_/A vssd1 vssd1 vccd1 vccd1 _3259_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6047_ _6749_/Q _5523_/X _6046_/X _6027_/X vssd1 vssd1 vccd1 vccd1 _6749_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6949_ _6949_/A _3247_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5280_ _6605_/Q _5282_/B vssd1 vssd1 vccd1 vccd1 _5281_/A sky130_fd_sc_hd__and2_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4300_ _4296_/X _4300_/B _4333_/A _4301_/A vssd1 vssd1 vccd1 vccd1 _4304_/B sky130_fd_sc_hd__and4b_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ _4231_/A _4231_/B vssd1 vssd1 vccd1 vccd1 _4232_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4162_ _4175_/A _4160_/X _4122_/B _4145_/Y vssd1 vssd1 vccd1 vccd1 _4162_/Y sky130_fd_sc_hd__a211oi_2
X_4093_ _4093_/A _4093_/B vssd1 vssd1 vccd1 vccd1 _4093_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4995_ _6548_/Q _4996_/B _4994_/X vssd1 vssd1 vccd1 vccd1 _6548_/D sky130_fd_sc_hd__o21ba_1
XFILLER_63_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6803_ _6809_/CLK _6803_/D vssd1 vssd1 vccd1 vccd1 _6803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6734_ _6809_/CLK _6734_/D vssd1 vssd1 vccd1 vccd1 _6734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3946_ _3944_/X _3946_/B vssd1 vssd1 vccd1 vccd1 _3947_/B sky130_fd_sc_hd__and2b_1
X_6665_ _6667_/CLK _6665_/D vssd1 vssd1 vccd1 vccd1 _6665_/Q sky130_fd_sc_hd__dfxtp_1
X_3877_ _5214_/C _4257_/B vssd1 vssd1 vccd1 vccd1 _3878_/A sky130_fd_sc_hd__and2_1
X_6596_ _6667_/CLK _6596_/D vssd1 vssd1 vccd1 vccd1 _6596_/Q sky130_fd_sc_hd__dfxtp_1
X_5616_ _6003_/A vssd1 vssd1 vccd1 vccd1 _5616_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5547_ _5542_/X _5525_/X _5505_/X _5546_/X vssd1 vssd1 vccd1 vccd1 _5547_/X sky130_fd_sc_hd__o211a_1
XFILLER_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5478_ _5490_/A _5478_/B vssd1 vssd1 vccd1 vccd1 _5479_/A sky130_fd_sc_hd__and2_1
X_4429_ _4429_/A _4450_/B _4429_/C vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__and3_1
XFILLER_59_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3800_ _3820_/A _3820_/B vssd1 vssd1 vccd1 vccd1 _3801_/B sky130_fd_sc_hd__xor2_2
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _4791_/A vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3731_ _3769_/A _3752_/B _3730_/X vssd1 vssd1 vccd1 vccd1 _3734_/A sky130_fd_sc_hd__o21bai_1
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3662_ _3706_/C _3662_/B vssd1 vssd1 vccd1 vccd1 _3663_/B sky130_fd_sc_hd__xnor2_1
X_6450_ _6789_/CLK _6450_/D vssd1 vssd1 vccd1 vccd1 _6450_/Q sky130_fd_sc_hd__dfxtp_1
X_5401_ _5401_/A vssd1 vssd1 vccd1 vccd1 _6642_/D sky130_fd_sc_hd__clkbuf_1
X_6381_ _6795_/CLK _6381_/D vssd1 vssd1 vccd1 vccd1 _6381_/Q sky130_fd_sc_hd__dfxtp_1
X_3593_ _3593_/A _3593_/B _3591_/Y vssd1 vssd1 vccd1 vccd1 _3594_/C sky130_fd_sc_hd__or3b_1
X_5332_ _5329_/Y _5335_/B _5331_/X vssd1 vssd1 vccd1 vccd1 _6621_/D sky130_fd_sc_hd__o21ai_1
X_5263_ _6597_/Q _5271_/B vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__and2_1
X_5194_ _6921_/A _5209_/B vssd1 vssd1 vccd1 vccd1 _5197_/B sky130_fd_sc_hd__or2_1
XFILLER_87_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4214_ _4225_/B _4214_/B vssd1 vssd1 vccd1 vccd1 _4216_/B sky130_fd_sc_hd__xor2_1
XFILLER_95_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4145_ _4145_/A _4145_/B vssd1 vssd1 vccd1 vccd1 _4145_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4076_ _6663_/Q _4153_/B _4076_/C _4114_/C vssd1 vssd1 vccd1 vccd1 _4079_/C sky130_fd_sc_hd__nand4_1
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6821__81 vssd1 vssd1 vccd1 vccd1 _6821__81/HI _6930_/A sky130_fd_sc_hd__conb_1
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4978_ _4978_/A vssd1 vssd1 vccd1 vccd1 _6543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6717_ _6799_/CLK _6717_/D vssd1 vssd1 vccd1 vccd1 _6717_/Q sky130_fd_sc_hd__dfxtp_1
X_3929_ _3930_/A _3930_/B vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__or2_1
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6648_ _6763_/CLK _6648_/D vssd1 vssd1 vccd1 vccd1 _6648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6579_ _6580_/CLK _6579_/D vssd1 vssd1 vccd1 vccd1 _6917_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _5935_/X _5948_/X _5949_/X _5687_/X vssd1 vssd1 vccd1 vccd1 _5950_/X sky130_fd_sc_hd__a211o_1
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4901_ _6520_/Q _4870_/A _4873_/A input48/X vssd1 vssd1 vccd1 vccd1 _6520_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5881_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5964_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4832_ _6431_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4833_/A sky130_fd_sc_hd__and2_1
XFILLER_60_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4763_ _6400_/Q _4767_/B vssd1 vssd1 vccd1 vccd1 _4764_/A sky130_fd_sc_hd__and2_1
XFILLER_119_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6502_ _6504_/CLK _6502_/D vssd1 vssd1 vccd1 vccd1 _6502_/Q sky130_fd_sc_hd__dfxtp_1
X_3714_ _3715_/A _3828_/A vssd1 vssd1 vccd1 vccd1 _3716_/B sky130_fd_sc_hd__nand2_1
X_4694_ _6361_/Q _4700_/B vssd1 vssd1 vccd1 vccd1 _4695_/A sky130_fd_sc_hd__and2_1
XFILLER_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6433_ _6795_/CLK _6433_/D vssd1 vssd1 vccd1 vccd1 _6433_/Q sky130_fd_sc_hd__dfxtp_1
X_3645_ _6653_/Q _3645_/B vssd1 vssd1 vccd1 vccd1 _3647_/A sky130_fd_sc_hd__and2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3576_ _3576_/A _3576_/B vssd1 vssd1 vccd1 vccd1 _3599_/A sky130_fd_sc_hd__xnor2_1
X_6364_ _6763_/CLK _6364_/D vssd1 vssd1 vccd1 vccd1 _6364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6295_ _6570_/CLK _6295_/D vssd1 vssd1 vccd1 vccd1 _6295_/Q sky130_fd_sc_hd__dfxtp_1
X_5315_ _3349_/X _5406_/A _5406_/B _3352_/X vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__a31o_1
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5246_ _5879_/A _5246_/B vssd1 vssd1 vccd1 vccd1 _6589_/D sky130_fd_sc_hd__nor2_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5177_ _5150_/X _5175_/X _5176_/X vssd1 vssd1 vccd1 vccd1 _5178_/C sky130_fd_sc_hd__a21o_1
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4128_ _4128_/A _4128_/B _4128_/C vssd1 vssd1 vccd1 vccd1 _4144_/B sky130_fd_sc_hd__nand3_2
XFILLER_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4059_ _4103_/C _4059_/B vssd1 vssd1 vccd1 vccd1 _4060_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3430_ _3789_/C vssd1 vssd1 vccd1 vccd1 _3758_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3361_ _6551_/Q _6550_/Q _4928_/A vssd1 vssd1 vccd1 vccd1 _3361_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5100_ _6136_/A vssd1 vssd1 vccd1 vccd1 _5100_/X sky130_fd_sc_hd__clkbuf_4
X_6080_ _6106_/A vssd1 vssd1 vccd1 vccd1 _6080_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3292_ _3292_/A vssd1 vssd1 vccd1 vccd1 _3292_/Y sky130_fd_sc_hd__inv_2
X_5031_ _5043_/A _5031_/B vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__or2_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6982_ _6982_/A _3286_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
X_5933_ _5999_/A vssd1 vssd1 vccd1 vccd1 _5933_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5864_ _6718_/Q _5850_/X _5861_/X _5863_/X vssd1 vssd1 vccd1 vccd1 _6718_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4815_ _6423_/Q _4823_/B vssd1 vssd1 vccd1 vccd1 _4816_/A sky130_fd_sc_hd__and2_1
X_5795_ _6479_/Q _5787_/X _5794_/X _5777_/X _5788_/X vssd1 vssd1 vccd1 vccd1 _5795_/X
+ sky130_fd_sc_hd__a221o_1
X_4746_ _5284_/A vssd1 vssd1 vccd1 vccd1 _4791_/A sky130_fd_sc_hd__clkbuf_4
X_4677_ _6346_/Q _4677_/B vssd1 vssd1 vccd1 vccd1 _4678_/A sky130_fd_sc_hd__and2_1
X_3628_ _3591_/A _3591_/B _3627_/Y vssd1 vssd1 vccd1 vccd1 _3629_/C sky130_fd_sc_hd__a21o_1
X_6416_ _6763_/CLK _6416_/D vssd1 vssd1 vccd1 vccd1 _6416_/Q sky130_fd_sc_hd__dfxtp_1
X_6347_ _6789_/CLK _6347_/D vssd1 vssd1 vccd1 vccd1 _6347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3559_ _3559_/A _3559_/B vssd1 vssd1 vccd1 vccd1 _3571_/B sky130_fd_sc_hd__xnor2_2
XFILLER_102_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6278_ _6268_/X _6277_/Y _6264_/X vssd1 vssd1 vccd1 vccd1 _6278_/Y sky130_fd_sc_hd__o21ai_1
X_5229_ _5229_/A _5229_/B _5229_/C vssd1 vssd1 vccd1 vccd1 _5230_/D sky130_fd_sc_hd__or3_1
XFILLER_76_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4600_ _4600_/A _4600_/B _4600_/C vssd1 vssd1 vccd1 vccd1 _4601_/B sky130_fd_sc_hd__nor3_1
XFILLER_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5580_ _6677_/Q _5551_/X _5576_/X _5579_/X _5540_/X vssd1 vssd1 vccd1 vccd1 _6677_/D
+ sky130_fd_sc_hd__o221a_1
X_4531_ _4531_/A _4531_/B _4531_/C vssd1 vssd1 vccd1 vccd1 _4535_/B sky130_fd_sc_hd__nand3_1
X_4462_ _4460_/X _4462_/B vssd1 vssd1 vccd1 vccd1 _4462_/X sky130_fd_sc_hd__and2b_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3413_ _5217_/C _6501_/Q _3427_/S vssd1 vssd1 vccd1 vccd1 _3414_/A sky130_fd_sc_hd__mux2_1
X_6201_ _6790_/Q _6194_/X _6200_/X _6190_/X vssd1 vssd1 vccd1 vccd1 _6790_/D sky130_fd_sc_hd__o211a_1
X_4393_ _4543_/A _4479_/B _4393_/C _4550_/C vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__nand4_2
XFILLER_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6132_ _6132_/A _6132_/B vssd1 vssd1 vccd1 vccd1 _6133_/A sky130_fd_sc_hd__and2_1
X_3344_ _6461_/Q _6460_/Q _6459_/Q _6458_/Q vssd1 vssd1 vccd1 vccd1 _3346_/B sky130_fd_sc_hd__or4_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3281_/A vssd1 vssd1 vccd1 vccd1 _3280_/A sky130_fd_sc_hd__buf_8
XFILLER_97_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6841__101 vssd1 vssd1 vccd1 vccd1 _6841__101/HI _6950_/A sky130_fd_sc_hd__conb_1
X_6063_ _6113_/A vssd1 vssd1 vccd1 vccd1 _6138_/S sky130_fd_sc_hd__clkbuf_4
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5169_/A vssd1 vssd1 vccd1 vccd1 _5014_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _6965_/A _3266_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
XFILLER_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5916_ _5906_/X _5913_/X _5914_/X _5915_/X vssd1 vssd1 vccd1 vccd1 _5916_/X sky130_fd_sc_hd__a211o_1
X_6896_ _6896_/A _3310_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__ebufn_8
XFILLER_22_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5847_ _5630_/X _5846_/X _5860_/S vssd1 vssd1 vccd1 vccd1 _5847_/X sky130_fd_sc_hd__mux2_1
X_5778_ _6636_/Q _5778_/B _6637_/Q vssd1 vssd1 vccd1 vccd1 _5865_/S sky130_fd_sc_hd__and3b_2
XFILLER_21_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4729_ _6385_/Q _4733_/B vssd1 vssd1 vccd1 vccd1 _4730_/A sky130_fd_sc_hd__and2_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6750_ _6799_/CLK _6750_/D vssd1 vssd1 vccd1 vccd1 _6750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5701_ _6690_/Q _5544_/X _5724_/S vssd1 vssd1 vccd1 vccd1 _5702_/B sky130_fd_sc_hd__mux2_1
X_3962_ _4058_/A _4268_/A vssd1 vssd1 vccd1 vccd1 _3963_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6681_ _6532_/Q _6681_/D vssd1 vssd1 vccd1 vccd1 _6681_/Q sky130_fd_sc_hd__dfxtp_1
X_3893_ _3992_/A vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5632_ _5632_/A vssd1 vssd1 vccd1 vccd1 _5670_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5563_ _5575_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _5563_/X sky130_fd_sc_hd__or2_1
X_4514_ _4514_/A _4553_/B _4514_/C vssd1 vssd1 vccd1 vccd1 _4557_/A sky130_fd_sc_hd__and3_1
X_5494_ _6084_/A _5494_/B vssd1 vssd1 vccd1 vccd1 _5495_/A sky130_fd_sc_hd__and2_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4445_ _4445_/A _4445_/B _4445_/C vssd1 vssd1 vccd1 vccd1 _4468_/C sky130_fd_sc_hd__nand3_1
X_4376_ _4404_/A _4376_/B vssd1 vssd1 vccd1 vccd1 _4390_/B sky130_fd_sc_hd__nor2_1
X_3327_ _3327_/A _3327_/B input5/X input4/X vssd1 vssd1 vccd1 vccd1 _3329_/C sky130_fd_sc_hd__or4_1
X_6115_ _6761_/Q _6106_/X _6114_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6116_/B sky130_fd_sc_hd__a22o_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3262_/A vssd1 vssd1 vccd1 vccd1 _3258_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6046_ _6029_/X _6044_/X _6045_/X vssd1 vssd1 vccd1 vccd1 _6046_/X sky130_fd_sc_hd__a21o_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3189_ _3193_/A vssd1 vssd1 vccd1 vccd1 _3189_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _6948_/A _3246_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4230_ _4242_/A _4241_/A _4230_/C _4230_/D vssd1 vssd1 vccd1 vccd1 _4231_/B sky130_fd_sc_hd__nand4_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4161_ _4122_/B _4145_/Y _4175_/A _4160_/X vssd1 vssd1 vccd1 vccd1 _4176_/B sky130_fd_sc_hd__o211a_1
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4092_ _4091_/A _4091_/B _4091_/C vssd1 vssd1 vccd1 vccd1 _4098_/C sky130_fd_sc_hd__a21o_1
XFILLER_83_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6802_ _6809_/CLK _6802_/D vssd1 vssd1 vccd1 vccd1 _6802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4994_ _6548_/Q _4993_/A _5017_/A _4993_/C _4385_/A vssd1 vssd1 vccd1 vccd1 _4994_/X
+ sky130_fd_sc_hd__a41o_1
X_6733_ _6799_/CLK _6733_/D vssd1 vssd1 vccd1 vccd1 _6733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3945_ _3944_/A _6350_/Q _4005_/D _3944_/B vssd1 vssd1 vccd1 vccd1 _3946_/B sky130_fd_sc_hd__a22o_1
X_6664_ _6667_/CLK _6664_/D vssd1 vssd1 vccd1 vccd1 _6664_/Q sky130_fd_sc_hd__dfxtp_1
X_5615_ _6487_/Q vssd1 vssd1 vccd1 vccd1 _6263_/A sky130_fd_sc_hd__buf_4
X_3876_ _3876_/A vssd1 vssd1 vccd1 vccd1 _6354_/D sky130_fd_sc_hd__clkbuf_1
X_6595_ _6667_/CLK _6595_/D vssd1 vssd1 vccd1 vccd1 _6595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5546_ _5575_/A _5546_/B vssd1 vssd1 vccd1 vccd1 _5546_/X sky130_fd_sc_hd__or2_1
XFILLER_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5477_ _6313_/Q _4499_/A _5483_/S vssd1 vssd1 vccd1 vccd1 _5478_/B sky130_fd_sc_hd__mux2_1
X_4428_ _4428_/A _4428_/B _4428_/C vssd1 vssd1 vccd1 vccd1 _4428_/Y sky130_fd_sc_hd__nand3_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4359_ _4388_/C _4359_/B vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6029_ _6029_/A vssd1 vssd1 vccd1 vccd1 _6029_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3730_ _3751_/A _3751_/B vssd1 vssd1 vccd1 vccd1 _3730_/X sky130_fd_sc_hd__xor2_1
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3661_ _3661_/A _3792_/B vssd1 vssd1 vccd1 vccd1 _3662_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5400_ _6642_/Q _5412_/B vssd1 vssd1 vccd1 vccd1 _5401_/A sky130_fd_sc_hd__and2_1
X_6380_ _6795_/CLK _6380_/D vssd1 vssd1 vccd1 vccd1 _6380_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3592_ _3593_/A _3593_/B _3591_/Y vssd1 vssd1 vccd1 vccd1 _3592_/X sky130_fd_sc_hd__o21ba_1
X_5331_ _5422_/A vssd1 vssd1 vccd1 vccd1 _5331_/X sky130_fd_sc_hd__buf_2
XFILLER_114_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5262_ _5273_/A vssd1 vssd1 vccd1 vccd1 _5271_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5193_ _5193_/A vssd1 vssd1 vccd1 vccd1 _5243_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4213_ _4192_/A _4192_/B _4212_/Y vssd1 vssd1 vccd1 vccd1 _4214_/B sky130_fd_sc_hd__a21boi_4
X_4144_ _4144_/A _4144_/B _4144_/C vssd1 vssd1 vccd1 vccd1 _4144_/Y sky130_fd_sc_hd__nand3_1
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4075_ _6663_/Q _4076_/C _6352_/Q _6662_/Q vssd1 vssd1 vccd1 vccd1 _4079_/B sky130_fd_sc_hd__a22o_1
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4977_ _6543_/Q _5249_/B vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__and2_1
X_6716_ _6799_/CLK _6716_/D vssd1 vssd1 vccd1 vccd1 _6716_/Q sky130_fd_sc_hd__dfxtp_1
X_3928_ _3928_/A _3928_/B vssd1 vssd1 vccd1 vccd1 _3930_/B sky130_fd_sc_hd__nor2_1
X_6647_ _6799_/CLK _6647_/D vssd1 vssd1 vccd1 vccd1 _6647_/Q sky130_fd_sc_hd__dfxtp_2
X_3859_ _3857_/X _3846_/X _3848_/Y _5001_/A vssd1 vssd1 vccd1 vccd1 _3860_/B sky130_fd_sc_hd__a31o_1
X_6578_ _6580_/CLK _6578_/D vssd1 vssd1 vccd1 vccd1 _6916_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5529_ _6447_/Q _5603_/B vssd1 vssd1 vccd1 vccd1 _5529_/X sky130_fd_sc_hd__and2_1
XFILLER_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4900_ _6519_/Q _4894_/X _4895_/X input46/X vssd1 vssd1 vccd1 vccd1 _6519_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5880_ _5880_/A _5880_/B vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__and2_2
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4831_ _4831_/A vssd1 vssd1 vccd1 vccd1 _6478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4762_ _4762_/A vssd1 vssd1 vccd1 vccd1 _6447_/D sky130_fd_sc_hd__clkbuf_1
X_3713_ _3674_/A _3676_/B _3673_/X vssd1 vssd1 vccd1 vccd1 _3828_/A sky130_fd_sc_hd__o21a_1
X_6501_ _6504_/CLK _6501_/D vssd1 vssd1 vccd1 vccd1 _6501_/Q sky130_fd_sc_hd__dfxtp_1
X_4693_ _4693_/A vssd1 vssd1 vccd1 vccd1 _6416_/D sky130_fd_sc_hd__clkbuf_1
X_6432_ _6795_/CLK _6432_/D vssd1 vssd1 vccd1 vccd1 _6432_/Q sky130_fd_sc_hd__dfxtp_1
X_3644_ _3789_/A _3759_/A _3681_/D _3644_/D vssd1 vssd1 vccd1 vccd1 _3647_/C sky130_fd_sc_hd__nand4_1
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6363_ _6763_/CLK _6363_/D vssd1 vssd1 vccd1 vccd1 _6363_/Q sky130_fd_sc_hd__dfxtp_1
X_3575_ _3616_/A _3808_/D vssd1 vssd1 vccd1 vccd1 _3576_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6294_ _6570_/CLK _6294_/D vssd1 vssd1 vccd1 vccd1 _6294_/Q sky130_fd_sc_hd__dfxtp_1
X_5314_ _6620_/Q vssd1 vssd1 vccd1 vccd1 _5502_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5245_ _6588_/Q _5242_/B _6589_/Q vssd1 vssd1 vccd1 vccd1 _5246_/B sky130_fd_sc_hd__a21oi_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5176_ _5176_/A vssd1 vssd1 vccd1 vccd1 _5176_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4127_ _4089_/A _4089_/C _4089_/B vssd1 vssd1 vccd1 vccd1 _4128_/C sky130_fd_sc_hd__a21bo_1
XFILLER_71_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4058_ _4058_/A _4058_/B vssd1 vssd1 vccd1 vccd1 _4059_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3360_ _6332_/Q vssd1 vssd1 vccd1 vccd1 _4928_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3292_/A vssd1 vssd1 vccd1 vccd1 _3291_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5030_ _6674_/Q _6706_/Q _6738_/Q _6770_/Q _5012_/X _5029_/X vssd1 vssd1 vccd1 vccd1
+ _5031_/B sky130_fd_sc_hd__mux4_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6981_ _6981_/A _3285_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
XFILLER_26_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5932_ _5906_/X _5930_/X _5931_/X _5915_/X vssd1 vssd1 vccd1 vccd1 _5932_/X sky130_fd_sc_hd__a211o_1
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5863_ _5999_/A vssd1 vssd1 vccd1 vccd1 _5863_/X sky130_fd_sc_hd__buf_2
X_4814_ _4847_/A vssd1 vssd1 vccd1 vccd1 _4823_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5794_ _5524_/X _5792_/X _5814_/S vssd1 vssd1 vccd1 vccd1 _5794_/X sky130_fd_sc_hd__mux2_1
X_4745_ _4745_/A vssd1 vssd1 vccd1 vccd1 _6440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4676_ _4676_/A vssd1 vssd1 vccd1 vccd1 _6409_/D sky130_fd_sc_hd__clkbuf_1
X_3627_ _3627_/A _3627_/B vssd1 vssd1 vccd1 vccd1 _3627_/Y sky130_fd_sc_hd__nor2_1
X_6415_ _6809_/CLK _6415_/D vssd1 vssd1 vccd1 vccd1 _6415_/Q sky130_fd_sc_hd__dfxtp_1
X_6346_ _6789_/CLK _6346_/D vssd1 vssd1 vccd1 vccd1 _6346_/Q sky130_fd_sc_hd__dfxtp_1
X_3558_ _3556_/X _3558_/B vssd1 vssd1 vccd1 vccd1 _3559_/B sky130_fd_sc_hd__and2b_1
XFILLER_103_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3489_ _6322_/Q _6526_/Q _3495_/S vssd1 vssd1 vccd1 vccd1 _3490_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6277_ _6277_/A _6283_/B vssd1 vssd1 vccd1 vccd1 _6277_/Y sky130_fd_sc_hd__nand2_1
X_5228_ _6606_/Q _6605_/Q _6603_/Q _6602_/Q vssd1 vssd1 vccd1 vccd1 _5229_/C sky130_fd_sc_hd__or4_1
XFILLER_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5159_ _5150_/X _5158_/X _5145_/X vssd1 vssd1 vccd1 vccd1 _5160_/C sky130_fd_sc_hd__a21o_1
XFILLER_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4530_ _4527_/Y _4528_/X _4493_/B _4493_/Y vssd1 vssd1 vccd1 vccd1 _4531_/C sky130_fd_sc_hd__o211ai_2
XFILLER_116_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4461_ _4416_/B _4420_/A _4458_/Y _4459_/X vssd1 vssd1 vccd1 vccd1 _4462_/B sky130_fd_sc_hd__a211o_1
X_3412_ _3516_/D vssd1 vssd1 vccd1 vccd1 _5217_/C sky130_fd_sc_hd__clkbuf_2
X_6200_ _6253_/A _6205_/B vssd1 vssd1 vccd1 vccd1 _6200_/X sky130_fd_sc_hd__or2_1
XFILLER_112_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4392_ _4368_/A _4510_/C _4550_/C _4368_/B vssd1 vssd1 vccd1 vccd1 _4396_/C sky130_fd_sc_hd__a22o_1
X_6131_ _6765_/Q _6106_/A _6130_/X _5406_/C vssd1 vssd1 vccd1 vccd1 _6132_/B sky130_fd_sc_hd__a22o_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _6457_/Q _6456_/Q _6455_/Q _6454_/Q vssd1 vssd1 vccd1 vccd1 _3346_/A sky130_fd_sc_hd__or4_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6062_ _6622_/Q _6224_/C _6062_/C vssd1 vssd1 vccd1 vccd1 _6113_/A sky130_fd_sc_hd__and3_2
X_6880__140 vssd1 vssd1 vccd1 vccd1 _6880__140/HI _6989_/A sky130_fd_sc_hd__conb_1
X_3274_ _3274_/A vssd1 vssd1 vccd1 vccd1 _3274_/Y sky130_fd_sc_hd__inv_2
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _6534_/Q vssd1 vssd1 vccd1 vccd1 _5169_/A sky130_fd_sc_hd__buf_4
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6964_ _6964_/A _3265_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
X_5915_ _5915_/A vssd1 vssd1 vccd1 vccd1 _5915_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6895_ _6895_/A _3183_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__ebufn_8
X_5846_ _6715_/Q _5633_/X _5859_/S vssd1 vssd1 vccd1 vccd1 _5846_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5777_ _5836_/A vssd1 vssd1 vccd1 vccd1 _5777_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4728_ _4728_/A vssd1 vssd1 vccd1 vccd1 _6432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4659_ _4659_/A vssd1 vssd1 vccd1 vccd1 _6401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6329_ _6799_/CLK _6329_/D vssd1 vssd1 vccd1 vccd1 _6329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6864__124 vssd1 vssd1 vccd1 vccd1 _6864__124/HI _6973_/A sky130_fd_sc_hd__conb_1
XFILLER_106_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ _4123_/A _3998_/C _3946_/B _3944_/X vssd1 vssd1 vccd1 vccd1 _3992_/C sky130_fd_sc_hd__a31o_1
XFILLER_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5700_ _5700_/A _6059_/A vssd1 vssd1 vccd1 vccd1 _5765_/A sky130_fd_sc_hd__nor2_2
X_6680_ _6532_/Q _6680_/D vssd1 vssd1 vccd1 vccd1 _6680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3892_ _4058_/A vssd1 vssd1 vccd1 vccd1 _3992_/A sky130_fd_sc_hd__clkbuf_2
X_5631_ _5631_/A vssd1 vssd1 vccd1 vccd1 _5631_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5562_ _6676_/Q _5561_/X _5562_/S vssd1 vssd1 vccd1 vccd1 _5563_/B sky130_fd_sc_hd__mux2_1
X_4513_ _4473_/A _4473_/B _4473_/C vssd1 vssd1 vccd1 vccd1 _4514_/C sky130_fd_sc_hd__a21bo_1
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5493_ _6318_/Q _4636_/A _5496_/S vssd1 vssd1 vccd1 vccd1 _5494_/B sky130_fd_sc_hd__mux2_1
XFILLER_7_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4444_ _4445_/B _4445_/C _4445_/A vssd1 vssd1 vccd1 vccd1 _4468_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4375_ _4597_/A _4373_/D _4369_/X _4371_/X vssd1 vssd1 vccd1 vccd1 _4376_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3326_ _3326_/A input3/X _3326_/C _3326_/D vssd1 vssd1 vccd1 vccd1 _3329_/B sky130_fd_sc_hd__or4_1
X_6114_ _6471_/Q _6107_/X _6096_/X _6113_/X _6487_/Q vssd1 vssd1 vccd1 vccd1 _6114_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6491_/Q _6023_/X _6249_/A _6031_/X vssd1 vssd1 vccd1 vccd1 _6045_/X sky130_fd_sc_hd__a31o_1
X_6828__88 vssd1 vssd1 vccd1 vccd1 _6828__88/HI _6937_/A sky130_fd_sc_hd__conb_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3281_/A vssd1 vssd1 vccd1 vccd1 _3262_/A sky130_fd_sc_hd__buf_12
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3193_/A sky130_fd_sc_hd__buf_2
XFILLER_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6947_ _6947_/A _3245_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5829_ _6711_/Q _5825_/X _5828_/X _5810_/X vssd1 vssd1 vccd1 vccd1 _6711_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6848__108 vssd1 vssd1 vccd1 vccd1 _6848__108/HI _6957_/A sky130_fd_sc_hd__conb_1
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4160_ _4160_/A _4160_/B _4160_/C vssd1 vssd1 vccd1 vccd1 _4160_/X sky130_fd_sc_hd__or3_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4091_ _4091_/A _4091_/B _4091_/C vssd1 vssd1 vccd1 vccd1 _4098_/B sky130_fd_sc_hd__nand3_2
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6801_ _6809_/CLK _6801_/D vssd1 vssd1 vccd1 vccd1 _6801_/Q sky130_fd_sc_hd__dfxtp_1
X_4993_ _4993_/A _5008_/C _4993_/C vssd1 vssd1 vccd1 vccd1 _4996_/B sky130_fd_sc_hd__and3_1
XFILLER_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6732_ _6799_/CLK _6732_/D vssd1 vssd1 vccd1 vccd1 _6732_/Q sky130_fd_sc_hd__dfxtp_1
X_3944_ _3944_/A _3944_/B _6350_/Q _4005_/D vssd1 vssd1 vccd1 vccd1 _3944_/X sky130_fd_sc_hd__and4_1
X_6663_ _6795_/CLK _6663_/D vssd1 vssd1 vccd1 vccd1 _6663_/Q sky130_fd_sc_hd__dfxtp_2
X_3875_ _5214_/D _4257_/B vssd1 vssd1 vccd1 vccd1 _3876_/A sky130_fd_sc_hd__and2_1
X_5614_ _5610_/X _5582_/X _5571_/X _5613_/X vssd1 vssd1 vccd1 vccd1 _5614_/X sky130_fd_sc_hd__o211a_1
X_6594_ _6667_/CLK _6594_/D vssd1 vssd1 vccd1 vccd1 _6594_/Q sky130_fd_sc_hd__dfxtp_1
X_5545_ _6674_/Q _5544_/X _5562_/S vssd1 vssd1 vccd1 vccd1 _5546_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5476_ _6112_/A vssd1 vssd1 vccd1 vccd1 _5490_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4427_ _4427_/A _4411_/B vssd1 vssd1 vccd1 vccd1 _4427_/X sky130_fd_sc_hd__or2b_1
X_4358_ _4451_/A _4388_/B vssd1 vssd1 vccd1 vccd1 _4359_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3309_ _3310_/A vssd1 vssd1 vccd1 vccd1 _3309_/Y sky130_fd_sc_hd__inv_2
X_4289_ _4400_/D vssd1 vssd1 vccd1 vccd1 _4296_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6028_ _6745_/Q _6011_/X _6025_/X _6027_/X vssd1 vssd1 vccd1 vccd1 _6745_/D sky130_fd_sc_hd__o211a_1
XFILLER_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3660_ _3660_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3706_/C sky130_fd_sc_hd__nand2_1
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3591_ _3591_/A _3591_/B vssd1 vssd1 vccd1 vccd1 _3591_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_114_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5330_ _5876_/B _5502_/B _5337_/B vssd1 vssd1 vccd1 vccd1 _5335_/B sky130_fd_sc_hd__and3_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5261_ _5261_/A vssd1 vssd1 vccd1 vccd1 _6596_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6554_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_114_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7000_ _7000_/A _3308_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
X_4212_ _4212_/A _4212_/B vssd1 vssd1 vccd1 vccd1 _4212_/Y sky130_fd_sc_hd__nand2_1
X_5192_ _5192_/A vssd1 vssd1 vccd1 vccd1 _6582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4143_ _4140_/Y _4141_/X _4142_/Y vssd1 vssd1 vccd1 vccd1 _6367_/D sky130_fd_sc_hd__a21oi_1
XFILLER_83_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4074_ _4074_/A _4074_/B _4074_/C vssd1 vssd1 vccd1 vccd1 _4074_/X sky130_fd_sc_hd__and3_1
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4976_ _5273_/A vssd1 vssd1 vccd1 vccd1 _5249_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6715_ _6799_/CLK _6715_/D vssd1 vssd1 vccd1 vccd1 _6715_/Q sky130_fd_sc_hd__dfxtp_1
X_3927_ _3927_/A _3927_/B vssd1 vssd1 vccd1 vccd1 _3930_/A sky130_fd_sc_hd__xnor2_1
XFILLER_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6646_ _6799_/CLK _6646_/D vssd1 vssd1 vccd1 vccd1 _6646_/Q sky130_fd_sc_hd__dfxtp_1
X_3858_ _3846_/X _3848_/Y _3857_/X vssd1 vssd1 vccd1 vccd1 _3860_/A sky130_fd_sc_hd__a21oi_2
XFILLER_118_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6577_ _6580_/CLK _6577_/D vssd1 vssd1 vccd1 vccd1 _6915_/A sky130_fd_sc_hd__dfxtp_1
X_3789_ _3789_/A _3789_/B _3789_/C _3789_/D vssd1 vssd1 vccd1 vccd1 _3813_/A sky130_fd_sc_hd__and4_1
X_5528_ _5668_/B vssd1 vssd1 vccd1 vccd1 _5603_/B sky130_fd_sc_hd__clkbuf_1
X_5459_ _6112_/A vssd1 vssd1 vccd1 vccd1 _5474_/A sky130_fd_sc_hd__buf_2
XFILLER_59_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4830_ _6430_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4831_/A sky130_fd_sc_hd__and2_1
XFILLER_61_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _6399_/Q _4767_/B vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__and2_1
XFILLER_119_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3712_ _3778_/A _3778_/B vssd1 vssd1 vccd1 vccd1 _3715_/A sky130_fd_sc_hd__or2_1
X_6500_ _6504_/CLK _6500_/D vssd1 vssd1 vccd1 vccd1 _6500_/Q sky130_fd_sc_hd__dfxtp_1
X_4692_ _6360_/Q _4700_/B vssd1 vssd1 vccd1 vccd1 _4693_/A sky130_fd_sc_hd__and2_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6431_ _6795_/CLK _6431_/D vssd1 vssd1 vccd1 vccd1 _6431_/Q sky130_fd_sc_hd__dfxtp_1
X_3643_ _6655_/Q vssd1 vssd1 vccd1 vccd1 _3789_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6362_ _6763_/CLK _6362_/D vssd1 vssd1 vccd1 vccd1 _6362_/Q sky130_fd_sc_hd__dfxtp_1
X_5313_ _5313_/A vssd1 vssd1 vccd1 vccd1 _6619_/D sky130_fd_sc_hd__clkbuf_1
X_3574_ _3596_/C _3574_/B vssd1 vssd1 vccd1 vccd1 _3576_/A sky130_fd_sc_hd__xnor2_1
X_6293_ _6584_/CLK _6293_/D vssd1 vssd1 vccd1 vccd1 _6293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5244_ _5244_/A vssd1 vssd1 vccd1 vccd1 _6588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5175_ _6697_/Q _6729_/Q _6761_/Q _6793_/Q _5157_/X _5169_/X vssd1 vssd1 vccd1 vccd1
+ _5175_/X sky130_fd_sc_hd__mux4_2
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _4160_/A _4146_/B _4124_/X vssd1 vssd1 vccd1 vccd1 _4128_/B sky130_fd_sc_hd__or3b_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _4057_/A _4057_/B vssd1 vssd1 vccd1 vccd1 _4103_/C sky130_fd_sc_hd__nand2_1
XFILLER_71_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4959_ _6537_/Q _4959_/B vssd1 vssd1 vccd1 vccd1 _4960_/A sky130_fd_sc_hd__and2_1
X_6629_ _6799_/CLK _6629_/D vssd1 vssd1 vccd1 vccd1 _6629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3290_ _3292_/A vssd1 vssd1 vccd1 vccd1 _3290_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6980_ _6980_/A _3284_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5931_ _6487_/Q _5931_/B _5943_/C vssd1 vssd1 vccd1 vccd1 _5931_/X sky130_fd_sc_hd__and3_1
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5862_ _6189_/A vssd1 vssd1 vccd1 vccd1 _5999_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4813_ _4813_/A vssd1 vssd1 vccd1 vccd1 _6470_/D sky130_fd_sc_hd__clkbuf_1
X_5793_ _5866_/S vssd1 vssd1 vccd1 vccd1 _5814_/S sky130_fd_sc_hd__clkbuf_2
X_4744_ _6392_/Q _4744_/B vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__and2_1
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4675_ _6345_/Q _4677_/B vssd1 vssd1 vccd1 vccd1 _4676_/A sky130_fd_sc_hd__and2_1
X_3626_ _3625_/B _3625_/C _3625_/A vssd1 vssd1 vccd1 vccd1 _3629_/B sky130_fd_sc_hd__o21ai_1
X_6414_ _6809_/CLK _6414_/D vssd1 vssd1 vccd1 vccd1 _6414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6345_ _6789_/CLK _6345_/D vssd1 vssd1 vccd1 vccd1 _6345_/Q sky130_fd_sc_hd__dfxtp_1
X_3557_ _3690_/B _3556_/C _3644_/D _3753_/A vssd1 vssd1 vccd1 vccd1 _3558_/B sky130_fd_sc_hd__a22o_1
X_6276_ _6811_/Q _6267_/X _6274_/Y _6275_/X vssd1 vssd1 vccd1 vccd1 _6811_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5227_ _6594_/Q _6593_/Q _6591_/Q _6590_/Q vssd1 vssd1 vccd1 vccd1 _5229_/B sky130_fd_sc_hd__or4_1
X_3488_ _3488_/A vssd1 vssd1 vccd1 vccd1 _6321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5158_ _6694_/Q _6726_/Q _6758_/Q _6790_/Q _5157_/X _5138_/X vssd1 vssd1 vccd1 vccd1
+ _5158_/X sky130_fd_sc_hd__mux4_2
X_5089_ _5081_/X _5085_/X _5087_/X _5088_/X vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__a31o_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4109_ _4168_/A _4168_/B vssd1 vssd1 vccd1 vccd1 _4109_/X sky130_fd_sc_hd__or2_1
XFILLER_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _4458_/Y _4459_/X _4416_/B _4420_/A vssd1 vssd1 vccd1 vccd1 _4460_/X sky130_fd_sc_hd__o211a_1
XFILLER_116_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4391_ _6377_/Q vssd1 vssd1 vccd1 vccd1 _4550_/C sky130_fd_sc_hd__clkbuf_2
X_3411_ _3556_/C vssd1 vssd1 vccd1 vccd1 _3516_/D sky130_fd_sc_hd__clkbuf_2
X_6130_ _6475_/Q _5919_/A _6070_/A _6113_/X _6491_/Q vssd1 vssd1 vccd1 vccd1 _6130_/X
+ sky130_fd_sc_hd__a32o_1
X_3342_ _6453_/Q _6452_/Q _6451_/Q _6450_/Q vssd1 vssd1 vccd1 vccd1 _3347_/A sky130_fd_sc_hd__or4_4
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3273_ _3274_/A vssd1 vssd1 vccd1 vccd1 _3273_/Y sky130_fd_sc_hd__inv_2
X_6061_ _6106_/A vssd1 vssd1 vccd1 vccd1 _6061_/X sky130_fd_sc_hd__clkbuf_4
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _6533_/Q vssd1 vssd1 vccd1 vccd1 _5012_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6963_ _6963_/A _3311_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
XFILLER_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5914_ _6484_/Q _5931_/B _5914_/C vssd1 vssd1 vccd1 vccd1 _5914_/X sky130_fd_sc_hd__and3_1
X_6894_ _6894_/A _3318_/A vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__ebufn_8
X_5845_ _6714_/Q _5825_/X _5844_/X _5838_/X vssd1 vssd1 vccd1 vccd1 _6714_/D sky130_fd_sc_hd__o211a_1
X_5776_ _6224_/A _5870_/B _6143_/B vssd1 vssd1 vccd1 vccd1 _5836_/A sky130_fd_sc_hd__or3_2
X_4727_ _6384_/Q _4733_/B vssd1 vssd1 vccd1 vccd1 _4728_/A sky130_fd_sc_hd__and2_1
X_4658_ _6337_/Q _4666_/B vssd1 vssd1 vccd1 vccd1 _4659_/A sky130_fd_sc_hd__and2_1
XFILLER_107_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3609_ _6297_/Q vssd1 vssd1 vccd1 vccd1 _3681_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4589_ _4593_/A _4593_/B vssd1 vssd1 vccd1 vccd1 _4590_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6328_ _6799_/CLK _6328_/D vssd1 vssd1 vccd1 vccd1 _6328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6259_ _6807_/Q _6247_/X _6258_/Y _6255_/X vssd1 vssd1 vccd1 vccd1 _6807_/D sky130_fd_sc_hd__o211a_1
XFILLER_76_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3960_ _6658_/Q vssd1 vssd1 vccd1 vccd1 _4123_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3891_ _6657_/Q vssd1 vssd1 vccd1 vccd1 _4058_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5630_ _6473_/Q vssd1 vssd1 vccd1 vccd1 _5630_/X sky130_fd_sc_hd__buf_2
X_5561_ _6450_/Q _5660_/B vssd1 vssd1 vccd1 vccd1 _5561_/X sky130_fd_sc_hd__and2_2
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4512_ _4547_/A _4512_/B _4512_/C _4553_/A vssd1 vssd1 vccd1 vccd1 _4553_/B sky130_fd_sc_hd__nand4_1
X_5492_ _6112_/A vssd1 vssd1 vccd1 vccd1 _6084_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_105_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4443_ _4487_/A _4487_/B vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__xor2_1
XFILLER_98_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4374_ _4547_/A vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__clkbuf_2
X_3325_ _3325_/A _3325_/B _3325_/C _3325_/D vssd1 vssd1 vccd1 vccd1 _3329_/A sky130_fd_sc_hd__or4_1
X_6113_ _6113_/A vssd1 vssd1 vccd1 vccd1 _6113_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ input1/X vssd1 vssd1 vccd1 vccd1 _3281_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6044_ _6749_/Q _5651_/X _6044_/S vssd1 vssd1 vccd1 vccd1 _6044_/X sky130_fd_sc_hd__mux2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _3187_/A vssd1 vssd1 vccd1 vccd1 _3187_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6946_ _6946_/A _3243_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5828_ _6485_/Q _5812_/X _5827_/X _5808_/X _5815_/X vssd1 vssd1 vccd1 vccd1 _5828_/X
+ sky130_fd_sc_hd__a221o_1
X_5759_ _6700_/Q _5755_/X _5758_/X _5739_/X vssd1 vssd1 vccd1 vccd1 _6700_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6887__147 vssd1 vssd1 vccd1 vccd1 _6887__147/HI _6996_/A sky130_fd_sc_hd__conb_1
XFILLER_108_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4090_ _4052_/A _4052_/C _4052_/B vssd1 vssd1 vccd1 vccd1 _4091_/C sky130_fd_sc_hd__a21bo_1
XFILLER_48_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6800_ _6809_/CLK _6800_/D vssd1 vssd1 vccd1 vccd1 _6800_/Q sky130_fd_sc_hd__dfxtp_1
X_4992_ _4992_/A vssd1 vssd1 vccd1 vccd1 _6547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6731_ _6799_/CLK _6731_/D vssd1 vssd1 vccd1 vccd1 _6731_/Q sky130_fd_sc_hd__dfxtp_1
X_3943_ _6351_/Q vssd1 vssd1 vccd1 vccd1 _4005_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6662_ _6795_/CLK _6662_/D vssd1 vssd1 vccd1 vccd1 _6662_/Q sky130_fd_sc_hd__dfxtp_1
X_3874_ _6189_/A vssd1 vssd1 vccd1 vccd1 _4257_/B sky130_fd_sc_hd__buf_2
X_5613_ _5624_/A _5613_/B vssd1 vssd1 vccd1 vccd1 _5613_/X sky130_fd_sc_hd__or2_1
X_6593_ _6667_/CLK _6593_/D vssd1 vssd1 vccd1 vccd1 _6593_/Q sky130_fd_sc_hd__dfxtp_1
X_5544_ _6448_/Q _5660_/B vssd1 vssd1 vccd1 vccd1 _5544_/X sky130_fd_sc_hd__and2_1
X_5475_ _5475_/A vssd1 vssd1 vccd1 vccd1 _6664_/D sky130_fd_sc_hd__clkbuf_1
X_4426_ _4426_/A _4410_/A vssd1 vssd1 vccd1 vccd1 _4426_/X sky130_fd_sc_hd__or2b_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4357_ _4519_/A _4393_/C _4339_/B _4337_/X vssd1 vssd1 vccd1 vccd1 _4388_/C sky130_fd_sc_hd__a31o_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3308_ _3310_/A vssd1 vssd1 vccd1 vccd1 _3308_/Y sky130_fd_sc_hd__inv_2
X_4288_ _6375_/Q vssd1 vssd1 vccd1 vccd1 _4400_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _3243_/A vssd1 vssd1 vccd1 vccd1 _3239_/Y sky130_fd_sc_hd__inv_2
X_6027_ _6178_/A vssd1 vssd1 vccd1 vccd1 _6027_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _6929_/A _3222_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_58_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3590_ _3627_/A _3627_/B vssd1 vssd1 vccd1 vccd1 _3591_/B sky130_fd_sc_hd__xor2_1
X_5260_ _6596_/Q _5260_/B vssd1 vssd1 vccd1 vccd1 _5261_/A sky130_fd_sc_hd__and2_1
XFILLER_114_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4211_ _4211_/A _4247_/A vssd1 vssd1 vccd1 vccd1 _4225_/B sky130_fd_sc_hd__nor2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5191_ _5191_/A _5191_/B _5191_/C vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__and3_1
XFILLER_95_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4142_ _4140_/Y _4141_/X _3781_/X vssd1 vssd1 vccd1 vccd1 _4142_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4073_ _4990_/A _4073_/B vssd1 vssd1 vccd1 vccd1 _6365_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4975_ _6542_/Q _4974_/A _4255_/X vssd1 vssd1 vccd1 vccd1 _6542_/D sky130_fd_sc_hd__o21a_1
XFILLER_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6714_ _6799_/CLK _6714_/D vssd1 vssd1 vccd1 vccd1 _6714_/Q sky130_fd_sc_hd__dfxtp_1
X_3926_ _3921_/Y _3936_/B _3925_/X vssd1 vssd1 vccd1 vccd1 _3927_/B sky130_fd_sc_hd__o21ai_1
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6645_ _6799_/CLK _6645_/D vssd1 vssd1 vccd1 vccd1 _6645_/Q sky130_fd_sc_hd__dfxtp_1
X_3857_ _3857_/A _3857_/B vssd1 vssd1 vccd1 vccd1 _3857_/X sky130_fd_sc_hd__or2_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6576_ _6580_/CLK _6576_/D vssd1 vssd1 vccd1 vccd1 _6914_/A sky130_fd_sc_hd__dfxtp_1
X_3788_ _3835_/A _3758_/B _3605_/B _3836_/A vssd1 vssd1 vccd1 vccd1 _3790_/A sky130_fd_sc_hd__a22oi_1
XFILLER_3_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5527_ _5632_/A vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5458_ _5458_/A vssd1 vssd1 vccd1 vccd1 _6112_/A sky130_fd_sc_hd__buf_2
X_4409_ _4451_/A _4595_/C vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__nand2_1
X_5389_ _5380_/X _5724_/S _5388_/Y _6067_/A vssd1 vssd1 vccd1 vccd1 _6636_/D sky130_fd_sc_hd__a211oi_1
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4760_ _4760_/A vssd1 vssd1 vccd1 vccd1 _6446_/D sky130_fd_sc_hd__clkbuf_1
X_3711_ _3708_/Y _3709_/X _3667_/X _3678_/Y vssd1 vssd1 vccd1 vccd1 _3778_/B sky130_fd_sc_hd__o211a_1
X_4691_ _4735_/A vssd1 vssd1 vccd1 vccd1 _4700_/B sky130_fd_sc_hd__clkbuf_1
X_6430_ _6795_/CLK _6430_/D vssd1 vssd1 vccd1 vccd1 _6430_/Q sky130_fd_sc_hd__dfxtp_1
X_3642_ _6654_/Q _3681_/D _3644_/D _6655_/Q vssd1 vssd1 vccd1 vccd1 _3647_/B sky130_fd_sc_hd__a22o_1
X_6361_ _6763_/CLK _6361_/D vssd1 vssd1 vccd1 vccd1 _6361_/Q sky130_fd_sc_hd__dfxtp_1
X_5312_ _6619_/Q _5346_/B vssd1 vssd1 vccd1 vccd1 _5313_/A sky130_fd_sc_hd__and2_1
X_3573_ _3661_/A _3722_/B vssd1 vssd1 vccd1 vccd1 _3574_/B sky130_fd_sc_hd__nand2_1
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6292_ _6584_/CLK _6292_/D vssd1 vssd1 vccd1 vccd1 _6292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5243_ _5243_/A _5243_/B _5243_/C vssd1 vssd1 vccd1 vccd1 _5244_/A sky130_fd_sc_hd__and3_1
X_5174_ _6918_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5178_/B sky130_fd_sc_hd__or2_1
XFILLER_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4125_ _4160_/A _4146_/B _4124_/X vssd1 vssd1 vccd1 vccd1 _4128_/A sky130_fd_sc_hd__o21bai_1
XFILLER_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4056_ _4056_/A _4101_/A vssd1 vssd1 vccd1 vccd1 _4060_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4958_ _4958_/A vssd1 vssd1 vccd1 vccd1 _6536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4889_ _6510_/Q _4887_/X _4888_/X input37/X vssd1 vssd1 vccd1 vccd1 _6510_/D sky130_fd_sc_hd__a22o_1
X_3909_ _3928_/B vssd1 vssd1 vccd1 vccd1 _3909_/Y sky130_fd_sc_hd__inv_2
X_6628_ _6799_/CLK _6628_/D vssd1 vssd1 vccd1 vccd1 _6628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6559_ _6562_/CLK _6559_/D vssd1 vssd1 vccd1 vccd1 _6897_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5930_ _5610_/X _5919_/X _5920_/X _5912_/X _6729_/Q vssd1 vssd1 vccd1 vccd1 _5930_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_53_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5861_ _6492_/Q _5840_/X _5860_/X _5836_/A _5843_/X vssd1 vssd1 vccd1 vccd1 _5861_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4812_ _6422_/Q _4812_/B vssd1 vssd1 vccd1 vccd1 _4813_/A sky130_fd_sc_hd__and2_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5792_ _6705_/Q _5529_/X _5813_/S vssd1 vssd1 vccd1 vccd1 _5792_/X sky130_fd_sc_hd__mux2_1
X_4743_ _4743_/A vssd1 vssd1 vccd1 vccd1 _6439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4674_ _4674_/A vssd1 vssd1 vccd1 vccd1 _6408_/D sky130_fd_sc_hd__clkbuf_1
X_6413_ _6789_/CLK _6413_/D vssd1 vssd1 vccd1 vccd1 _6413_/Q sky130_fd_sc_hd__dfxtp_1
X_3625_ _3625_/A _3625_/B _3625_/C vssd1 vssd1 vccd1 vccd1 _3629_/A sky130_fd_sc_hd__or3_1
X_6344_ _6789_/CLK _6344_/D vssd1 vssd1 vccd1 vccd1 _6344_/Q sky130_fd_sc_hd__dfxtp_1
X_3556_ _3753_/A _3690_/B _3556_/C _3644_/D vssd1 vssd1 vccd1 vccd1 _3556_/X sky130_fd_sc_hd__and4_1
XFILLER_115_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6275_ _6275_/A vssd1 vssd1 vccd1 vccd1 _6275_/X sky130_fd_sc_hd__clkbuf_2
X_5226_ _6601_/Q _6598_/Q _6597_/Q _6596_/Q vssd1 vssd1 vccd1 vccd1 _5229_/A sky130_fd_sc_hd__or4_1
X_3487_ _6321_/Q _6525_/Q _3495_/S vssd1 vssd1 vccd1 vccd1 _3488_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5157_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5088_ _5088_/A vssd1 vssd1 vccd1 vccd1 _5088_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4108_ _4105_/X _4106_/Y _4065_/B _4065_/Y vssd1 vssd1 vccd1 vccd1 _4168_/B sky130_fd_sc_hd__a211oi_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4039_ _4153_/A _4180_/B _4039_/C _4039_/D vssd1 vssd1 vccd1 vccd1 _4042_/C sky130_fd_sc_hd__nand4_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4390_ _4390_/A _4390_/B vssd1 vssd1 vccd1 vccd1 _4414_/A sky130_fd_sc_hd__nand2_1
X_3410_ _6297_/Q vssd1 vssd1 vccd1 vccd1 _3556_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3341_ _6331_/Q _3336_/X _3340_/X vssd1 vssd1 vccd1 vccd1 _6331_/D sky130_fd_sc_hd__o21a_1
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _3274_/A vssd1 vssd1 vccd1 vccd1 _3272_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6060_ _6058_/Y _6059_/X _5518_/A vssd1 vssd1 vccd1 vccd1 _6106_/A sky130_fd_sc_hd__a21o_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5011_ _5081_/A vssd1 vssd1 vccd1 vccd1 _5011_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6962_ _6962_/A _3264_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
X_5913_ _5581_/X _5889_/X _5891_/X _5912_/X _6726_/Q vssd1 vssd1 vccd1 vccd1 _5913_/X
+ sky130_fd_sc_hd__a32o_1
X_6893_ _6893_/A _3313_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__ebufn_8
X_5844_ _6488_/Q _5840_/X _5842_/X _5836_/X _5843_/X vssd1 vssd1 vccd1 vccd1 _5844_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5775_ _6620_/Q _5775_/B _5880_/A vssd1 vssd1 vccd1 vccd1 _6143_/B sky130_fd_sc_hd__or3b_4
X_4726_ _4726_/A vssd1 vssd1 vccd1 vccd1 _6431_/D sky130_fd_sc_hd__clkbuf_1
X_4657_ _4679_/A vssd1 vssd1 vccd1 vccd1 _4666_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3608_ _6654_/Q vssd1 vssd1 vccd1 vccd1 _3759_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6327_ _6528_/CLK _6327_/D vssd1 vssd1 vccd1 vccd1 _6327_/Q sky130_fd_sc_hd__dfxtp_1
X_4588_ _4588_/A _4588_/B vssd1 vssd1 vccd1 vccd1 _4593_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3539_ _3539_/A _3539_/B vssd1 vssd1 vccd1 vccd1 _3541_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6258_ _6248_/X _6257_/Y _6244_/X vssd1 vssd1 vccd1 vccd1 _6258_/Y sky130_fd_sc_hd__o21ai_1
X_5209_ _6924_/A _5209_/B vssd1 vssd1 vccd1 vccd1 _5212_/B sky130_fd_sc_hd__or2_1
X_6189_ _6189_/A vssd1 vssd1 vccd1 vccd1 _6255_/A sky130_fd_sc_hd__buf_2
XFILLER_123_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3890_ _3890_/A vssd1 vssd1 vccd1 vccd1 _6358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _6466_/Q vssd1 vssd1 vccd1 vccd1 _5560_/X sky130_fd_sc_hd__clkbuf_4
X_4511_ _6669_/Q _4576_/C _4512_/C _4553_/A vssd1 vssd1 vccd1 vccd1 _4514_/A sky130_fd_sc_hd__a22o_1
X_5491_ _5491_/A vssd1 vssd1 vccd1 vccd1 _6669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4442_ _4442_/A _4442_/B vssd1 vssd1 vccd1 vccd1 _4487_/B sky130_fd_sc_hd__or2_1
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4373_ _4369_/X _4371_/X _4547_/A _4373_/D vssd1 vssd1 vccd1 vccd1 _4404_/A sky130_fd_sc_hd__and4bb_1
X_3324_ _4941_/C _5008_/A _3324_/C _6892_/A vssd1 vssd1 vccd1 vccd1 _4993_/A sky130_fd_sc_hd__and4_1
X_6112_ _6112_/A vssd1 vssd1 vccd1 vccd1 _6132_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3255_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6043_ _6748_/Q _5523_/X _6042_/X _6027_/X vssd1 vssd1 vccd1 vccd1 _6748_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3187_/A vssd1 vssd1 vccd1 vccd1 _3186_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6945_ _6945_/A _3242_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5827_ _5593_/X _5826_/X _5842_/S vssd1 vssd1 vccd1 vccd1 _5827_/X sky130_fd_sc_hd__mux2_1
X_5758_ _6277_/A _5734_/X _5735_/X _5757_/X _5743_/X vssd1 vssd1 vccd1 vccd1 _5758_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4709_ _6368_/Q _4711_/B vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__and2_1
X_5689_ _6189_/A vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6819__79 vssd1 vssd1 vccd1 vccd1 _6819__79/HI _6928_/A sky130_fd_sc_hd__conb_1
XFILLER_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6870__130 vssd1 vssd1 vccd1 vccd1 _6870__130/HI _6979_/A sky130_fd_sc_hd__conb_1
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6833__93 vssd1 vssd1 vccd1 vccd1 _6833__93/HI _6942_/A sky130_fd_sc_hd__conb_1
XFILLER_76_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4991_ _6547_/Q _5249_/B vssd1 vssd1 vccd1 vccd1 _4992_/A sky130_fd_sc_hd__and2_1
X_6730_ _6799_/CLK _6730_/D vssd1 vssd1 vccd1 vccd1 _6730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _6660_/Q vssd1 vssd1 vccd1 vccd1 _3944_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6661_ _6795_/CLK _6661_/D vssd1 vssd1 vccd1 vccd1 _6661_/Q sky130_fd_sc_hd__dfxtp_2
X_3873_ _4259_/A vssd1 vssd1 vccd1 vccd1 _6189_/A sky130_fd_sc_hd__buf_2
X_6592_ _6667_/CLK _6592_/D vssd1 vssd1 vccd1 vccd1 _6592_/Q sky130_fd_sc_hd__dfxtp_1
X_5612_ _6681_/Q _5611_/X _5612_/S vssd1 vssd1 vccd1 vccd1 _5613_/B sky130_fd_sc_hd__mux2_1
X_5543_ _5668_/B vssd1 vssd1 vccd1 vccd1 _5660_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_117_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5474_ _5474_/A _5474_/B vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__and2_1
X_4425_ _4425_/A vssd1 vssd1 vccd1 vccd1 _6388_/D sky130_fd_sc_hd__clkbuf_1
X_4356_ _6666_/Q vssd1 vssd1 vccd1 vccd1 _4519_/A sky130_fd_sc_hd__clkbuf_2
X_3307_ _3310_/A vssd1 vssd1 vccd1 vccd1 _3307_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4287_ _4296_/A vssd1 vssd1 vccd1 vccd1 _4499_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _3250_/A vssd1 vssd1 vccd1 vccd1 _3243_/A sky130_fd_sc_hd__buf_12
XFILLER_104_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6026_ _6189_/A vssd1 vssd1 vccd1 vccd1 _6178_/A sky130_fd_sc_hd__buf_4
XFILLER_100_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6854__114 vssd1 vssd1 vccd1 vccd1 _6854__114/HI _6963_/A sky130_fd_sc_hd__conb_1
X_6928_ _6928_/A _3221_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4210_ _4210_/A _4210_/B vssd1 vssd1 vccd1 vccd1 _4247_/A sky130_fd_sc_hd__nor2_1
X_5190_ _5181_/X _5189_/X _5176_/X vssd1 vssd1 vccd1 vccd1 _5191_/C sky130_fd_sc_hd__a21o_1
X_4141_ _4109_/X _4220_/A _4168_/A vssd1 vssd1 vccd1 vccd1 _4141_/X sky130_fd_sc_hd__o21ba_1
XFILLER_110_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4072_ _4072_/A _4072_/B vssd1 vssd1 vccd1 vccd1 _4073_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4974_ _4974_/A _4974_/B vssd1 vssd1 vccd1 vccd1 _6541_/D sky130_fd_sc_hd__nor2_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3925_ _4058_/A _4264_/A _4266_/A _6656_/Q vssd1 vssd1 vccd1 vccd1 _3925_/X sky130_fd_sc_hd__a22o_1
X_6713_ _6532_/Q _6713_/D vssd1 vssd1 vccd1 vccd1 _6713_/Q sky130_fd_sc_hd__dfxtp_1
X_6644_ _6799_/CLK _6644_/D vssd1 vssd1 vccd1 vccd1 _6644_/Q sky130_fd_sc_hd__dfxtp_1
X_3856_ _3855_/A _3855_/B _3855_/C vssd1 vssd1 vccd1 vccd1 _3857_/B sky130_fd_sc_hd__a21oi_1
XFILLER_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6575_ _6580_/CLK _6575_/D vssd1 vssd1 vccd1 vccd1 _6913_/A sky130_fd_sc_hd__dfxtp_1
X_3787_ _3787_/A _3810_/B vssd1 vssd1 vccd1 vccd1 _3796_/A sky130_fd_sc_hd__nand2_1
X_5526_ _5873_/A _5700_/A vssd1 vssd1 vccd1 vccd1 _5632_/A sky130_fd_sc_hd__nor2_2
XFILLER_105_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5457_ _5457_/A vssd1 vssd1 vccd1 vccd1 _6659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4408_ _4477_/A _4371_/B _4371_/D _4368_/X vssd1 vssd1 vccd1 vccd1 _4410_/A sky130_fd_sc_hd__a31o_1
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5388_ _6011_/A _5778_/B _6636_/Q vssd1 vssd1 vccd1 vccd1 _5388_/Y sky130_fd_sc_hd__a21oi_1
X_4339_ _4337_/X _4339_/B vssd1 vssd1 vccd1 vccd1 _4340_/B sky130_fd_sc_hd__and2b_1
XFILLER_75_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6009_ _6001_/X _6007_/X _6008_/X vssd1 vssd1 vccd1 vccd1 _6009_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _3667_/X _3678_/Y _3708_/Y _3709_/X vssd1 vssd1 vccd1 vccd1 _3778_/A sky130_fd_sc_hd__a211oi_1
XFILLER_81_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4690_ _5458_/A vssd1 vssd1 vccd1 vccd1 _4735_/A sky130_fd_sc_hd__buf_2
X_3641_ _3641_/A _3660_/B _3641_/C vssd1 vssd1 vccd1 vccd1 _3679_/A sky130_fd_sc_hd__and3_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3572_ _3729_/A _3720_/D _3558_/B _3556_/X vssd1 vssd1 vccd1 vccd1 _3596_/C sky130_fd_sc_hd__a31o_1
X_6360_ _6763_/CLK _6360_/D vssd1 vssd1 vccd1 vccd1 _6360_/Q sky130_fd_sc_hd__dfxtp_1
X_5311_ _5311_/A vssd1 vssd1 vccd1 vccd1 _6618_/D sky130_fd_sc_hd__clkbuf_1
X_6291_ _6584_/CLK _6291_/D vssd1 vssd1 vccd1 vccd1 _6291_/Q sky130_fd_sc_hd__dfxtp_1
X_5242_ _6588_/Q _5242_/B vssd1 vssd1 vccd1 vccd1 _5243_/C sky130_fd_sc_hd__nand2_1
X_5173_ _5173_/A vssd1 vssd1 vccd1 vccd1 _6579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4124_ _4145_/A _4145_/B vssd1 vssd1 vccd1 vccd1 _4124_/X sky130_fd_sc_hd__xor2_1
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XFILLER_96_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4055_ _6357_/Q vssd1 vssd1 vccd1 vccd1 _4101_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4957_ _6536_/Q _4959_/B vssd1 vssd1 vccd1 vccd1 _4958_/A sky130_fd_sc_hd__and2_1
XFILLER_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4888_ _4895_/A vssd1 vssd1 vccd1 vccd1 _4888_/X sky130_fd_sc_hd__clkbuf_2
X_3908_ _3928_/A _3979_/D _3941_/A _3908_/D vssd1 vssd1 vccd1 vccd1 _3928_/B sky130_fd_sc_hd__and4b_1
X_6627_ _6532_/Q _6627_/D vssd1 vssd1 vccd1 vccd1 _6627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3839_ _3839_/A _3839_/B vssd1 vssd1 vccd1 vccd1 _3840_/B sky130_fd_sc_hd__nand2_1
X_6558_ _6558_/CLK _6558_/D vssd1 vssd1 vccd1 vccd1 _6896_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5509_ _6640_/Q _6639_/Q _6638_/Q _5509_/D vssd1 vssd1 vccd1 vccd1 _5510_/C sky130_fd_sc_hd__or4_2
X_6489_ _6795_/CLK _6489_/D vssd1 vssd1 vccd1 vccd1 _6489_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5860_ _5659_/X _5859_/X _5860_/S vssd1 vssd1 vccd1 vccd1 _5860_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4811_ _4811_/A vssd1 vssd1 vccd1 vccd1 _6469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5791_ _5865_/S vssd1 vssd1 vccd1 vccd1 _5813_/S sky130_fd_sc_hd__clkbuf_2
X_4742_ _6391_/Q _4744_/B vssd1 vssd1 vccd1 vccd1 _4743_/A sky130_fd_sc_hd__and2_1
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4673_ _6344_/Q _4677_/B vssd1 vssd1 vccd1 vccd1 _4674_/A sky130_fd_sc_hd__and2_1
X_3624_ _3671_/B _3671_/C _3671_/A vssd1 vssd1 vccd1 vccd1 _3625_/C sky130_fd_sc_hd__o21a_1
X_6412_ _6789_/CLK _6412_/D vssd1 vssd1 vccd1 vccd1 _6412_/Q sky130_fd_sc_hd__dfxtp_1
X_6343_ _6789_/CLK _6343_/D vssd1 vssd1 vccd1 vccd1 _6343_/Q sky130_fd_sc_hd__dfxtp_1
X_3555_ _6296_/Q vssd1 vssd1 vccd1 vccd1 _3644_/D sky130_fd_sc_hd__clkbuf_2
X_3486_ _3486_/A vssd1 vssd1 vccd1 vccd1 _3495_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6274_ _6268_/X _6273_/Y _6264_/X vssd1 vssd1 vccd1 vccd1 _6274_/Y sky130_fd_sc_hd__o21ai_1
X_5225_ _6614_/Q _6613_/Q _6612_/Q _6609_/Q vssd1 vssd1 vccd1 vccd1 _5230_/C sky130_fd_sc_hd__or4_1
XFILLER_69_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5156_ _6915_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5160_/B sky130_fd_sc_hd__or2_1
XFILLER_84_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5087_ _6810_/Q _5109_/B vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__or2_1
XFILLER_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4107_ _4065_/B _4065_/Y _4105_/X _4106_/Y vssd1 vssd1 vccd1 vccd1 _4168_/A sky130_fd_sc_hd__o211a_1
X_4038_ _4153_/A _6350_/Q _4005_/D _4180_/B vssd1 vssd1 vccd1 vccd1 _4042_/B sky130_fd_sc_hd__a22o_1
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _6738_/Q _5984_/X _5988_/X _5959_/X vssd1 vssd1 vccd1 vccd1 _6738_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_3340_ _5422_/A vssd1 vssd1 vccd1 vccd1 _3340_/X sky130_fd_sc_hd__buf_4
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3274_/A vssd1 vssd1 vccd1 vccd1 _3271_/Y sky130_fd_sc_hd__inv_2
X_5010_ _6554_/Q _6330_/Q _4255_/X vssd1 vssd1 vccd1 vccd1 _6554_/D sky130_fd_sc_hd__o21a_1
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6961_ _6961_/A _3262_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
X_6892_ _6892_/A _3309_/Y vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__ebufn_8
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5912_ _5941_/A vssd1 vssd1 vccd1 vccd1 _5912_/X sky130_fd_sc_hd__clkbuf_2
X_5843_ _5843_/A vssd1 vssd1 vccd1 vccd1 _5843_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5774_ _6703_/Q _5755_/X _5772_/X _5773_/X vssd1 vssd1 vccd1 vccd1 _6703_/D sky130_fd_sc_hd__o211a_1
X_4725_ _6383_/Q _4733_/B vssd1 vssd1 vccd1 vccd1 _4726_/A sky130_fd_sc_hd__and2_1
X_4656_ _4656_/A vssd1 vssd1 vccd1 vccd1 _6400_/D sky130_fd_sc_hd__clkbuf_1
X_4587_ _4607_/A _4607_/B vssd1 vssd1 vccd1 vccd1 _4588_/B sky130_fd_sc_hd__xor2_1
X_3607_ _3757_/A _3556_/C _3578_/B _3789_/B vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__a22oi_1
XFILLER_107_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6326_ _6531_/CLK _6326_/D vssd1 vssd1 vccd1 vccd1 _6326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3538_ _3538_/A _3538_/B vssd1 vssd1 vccd1 vccd1 _3541_/A sky130_fd_sc_hd__xnor2_1
XFILLER_115_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3469_ _6313_/Q _6517_/Q _3473_/S vssd1 vssd1 vccd1 vccd1 _3470_/A sky130_fd_sc_hd__mux2_1
X_6257_ _6257_/A _6263_/B vssd1 vssd1 vccd1 vccd1 _6257_/Y sky130_fd_sc_hd__nand2_1
X_5208_ _5208_/A vssd1 vssd1 vccd1 vccd1 _6585_/D sky130_fd_sc_hd__clkbuf_1
X_6188_ _6237_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _6188_/X sky130_fd_sc_hd__or2_1
XFILLER_123_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5139_ _6691_/Q _6723_/Q _6755_/Q _6787_/Q _5126_/X _5138_/X vssd1 vssd1 vccd1 vccd1
+ _5139_/X sky130_fd_sc_hd__mux4_2
XFILLER_57_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4510_ _4576_/A _4510_/B _4510_/C _4550_/C vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__nand4_1
X_5490_ _5490_/A _5490_/B vssd1 vssd1 vccd1 vccd1 _5491_/A sky130_fd_sc_hd__and2_1
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4441_ _4517_/A _4517_/B _6377_/Q _6378_/Q vssd1 vssd1 vccd1 vccd1 _4442_/B sky130_fd_sc_hd__and4_1
X_4372_ _6669_/Q vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__clkbuf_2
X_6111_ _6111_/A vssd1 vssd1 vccd1 vccd1 _6760_/D sky130_fd_sc_hd__clkbuf_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _6547_/Q _3323_/B vssd1 vssd1 vccd1 vccd1 _4980_/B sky130_fd_sc_hd__nor2_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6042_ _6029_/X _6039_/X _6041_/X vssd1 vssd1 vccd1 vccd1 _6042_/X sky130_fd_sc_hd__a21o_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3254_/Y sky130_fd_sc_hd__inv_2
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3185_ _3187_/A vssd1 vssd1 vccd1 vccd1 _3185_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6944_ _6944_/A _3241_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5826_ _6711_/Q _5594_/X _5841_/S vssd1 vssd1 vccd1 vccd1 _5826_/X sky130_fd_sc_hd__mux2_1
X_5757_ _5642_/X _5756_/X _5757_/S vssd1 vssd1 vccd1 vccd1 _5757_/X sky130_fd_sc_hd__mux2_1
X_4708_ _4708_/A vssd1 vssd1 vccd1 vccd1 _6423_/D sky130_fd_sc_hd__clkbuf_1
X_5688_ _6229_/A _5678_/X _5680_/X _5686_/X _5687_/X vssd1 vssd1 vccd1 vccd1 _5688_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4639_ _4627_/A _4626_/A _4626_/B _4638_/X vssd1 vssd1 vccd1 vccd1 _4640_/B sky130_fd_sc_hd__a31o_1
XFILLER_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6309_ _6522_/CLK _6309_/D vssd1 vssd1 vccd1 vccd1 _6309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4990_ _4990_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _6546_/D sky130_fd_sc_hd__nor2_1
XFILLER_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3941_ _3941_/A _4264_/A vssd1 vssd1 vccd1 vccd1 _3947_/A sky130_fd_sc_hd__nand2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6660_ _6795_/CLK _6660_/D vssd1 vssd1 vccd1 vccd1 _6660_/Q sky130_fd_sc_hd__dfxtp_1
X_3872_ _3872_/A vssd1 vssd1 vccd1 vccd1 _6353_/D sky130_fd_sc_hd__clkbuf_1
X_6591_ _6667_/CLK _6591_/D vssd1 vssd1 vccd1 vccd1 _6591_/Q sky130_fd_sc_hd__dfxtp_1
X_5611_ _6455_/Q _5652_/B vssd1 vssd1 vccd1 vccd1 _5611_/X sky130_fd_sc_hd__and2_2
X_5542_ _6464_/Q vssd1 vssd1 vccd1 vccd1 _5542_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5473_ _6312_/Q _4283_/A _5483_/S vssd1 vssd1 vccd1 vccd1 _5474_/B sky130_fd_sc_hd__mux2_1
X_4424_ _5129_/A _4424_/B _4463_/B vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__and3_1
XFILLER_113_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4355_ _4449_/A _4388_/B _4332_/A _4354_/X vssd1 vssd1 vccd1 vccd1 _4379_/A sky130_fd_sc_hd__a31o_1
XFILLER_86_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3306_ _3310_/A vssd1 vssd1 vccd1 vccd1 _3306_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4286_ _4451_/A vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6025_ _6001_/X _6022_/X _6024_/X vssd1 vssd1 vccd1 vccd1 _6025_/X sky130_fd_sc_hd__a21o_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3237_/A vssd1 vssd1 vccd1 vccd1 _3237_/Y sky130_fd_sc_hd__inv_2
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6927_ _6927_/A _3220_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_42_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5809_ _6482_/Q _5787_/X _5807_/X _5808_/X _5788_/X vssd1 vssd1 vccd1 vccd1 _5809_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6789_ _6789_/CLK _6789_/D vssd1 vssd1 vccd1 vccd1 _6789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4140_ _4140_/A _4140_/B vssd1 vssd1 vccd1 vccd1 _4140_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4071_ _3986_/X _4028_/B _4026_/X vssd1 vssd1 vccd1 vccd1 _4072_/B sky130_fd_sc_hd__a21oi_1
XFILLER_49_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6877__137 vssd1 vssd1 vccd1 vccd1 _6877__137/HI _6986_/A sky130_fd_sc_hd__conb_1
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _6541_/Q _4972_/B _4931_/X vssd1 vssd1 vccd1 vccd1 _4974_/B sky130_fd_sc_hd__o21ai_1
XFILLER_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3924_ _4058_/A _4266_/A vssd1 vssd1 vccd1 vccd1 _3936_/B sky130_fd_sc_hd__nand2_1
X_6712_ _6532_/Q _6712_/D vssd1 vssd1 vccd1 vccd1 _6712_/Q sky130_fd_sc_hd__dfxtp_1
X_6643_ _6667_/CLK _6643_/D vssd1 vssd1 vccd1 vccd1 _6643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3855_ _3855_/A _3855_/B _3855_/C vssd1 vssd1 vccd1 vccd1 _3857_/A sky130_fd_sc_hd__and3_1
XFILLER_118_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6574_ _6580_/CLK _6574_/D vssd1 vssd1 vccd1 vccd1 _6912_/A sky130_fd_sc_hd__dfxtp_1
X_3786_ _3786_/A _3786_/B vssd1 vssd1 vccd1 vccd1 _3806_/A sky130_fd_sc_hd__nor2_1
X_5525_ _5631_/A vssd1 vssd1 vccd1 vccd1 _5525_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5456_ _5456_/A _5456_/B vssd1 vssd1 vccd1 vccd1 _5457_/A sky130_fd_sc_hd__and2_1
X_4407_ _4407_/A _4579_/B vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5387_ _5770_/S vssd1 vssd1 vccd1 vccd1 _5724_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4338_ _4368_/A _4433_/C _4433_/D _4368_/B vssd1 vssd1 vccd1 vccd1 _4339_/B sky130_fd_sc_hd__a22o_1
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4269_ _4269_/A vssd1 vssd1 vccd1 vccd1 _6378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6008_ _6484_/Q _5996_/X _5986_/X _6003_/X vssd1 vssd1 vccd1 vccd1 _6008_/X sky130_fd_sc_hd__a31o_1
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3640_ _3671_/C vssd1 vssd1 vccd1 vccd1 _3640_/Y sky130_fd_sc_hd__inv_2
X_3571_ _3571_/A _3571_/B vssd1 vssd1 vccd1 vccd1 _3627_/A sky130_fd_sc_hd__nand2_1
X_6290_ _6584_/CLK _6290_/D vssd1 vssd1 vccd1 vccd1 _6290_/Q sky130_fd_sc_hd__dfxtp_1
X_5310_ _6618_/Q _5346_/B vssd1 vssd1 vccd1 vccd1 _5311_/A sky130_fd_sc_hd__and2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5241_ _6588_/Q _5242_/B vssd1 vssd1 vccd1 vccd1 _5243_/B sky130_fd_sc_hd__or2_1
XFILLER_123_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5172_ _5191_/A _5172_/B _5172_/C vssd1 vssd1 vccd1 vccd1 _5173_/A sky130_fd_sc_hd__and3_1
XFILLER_110_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4123_ _4123_/A _6357_/Q vssd1 vssd1 vccd1 vccd1 _4145_/B sky130_fd_sc_hd__nand2_1
Xinput2 wb_rst_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
XFILLER_110_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4054_ _4074_/B _4074_/C _4074_/A vssd1 vssd1 vccd1 vccd1 _4062_/C sky130_fd_sc_hd__a21o_1
XFILLER_71_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4956_ _5043_/A _4950_/X _4255_/X vssd1 vssd1 vccd1 vccd1 _6535_/D sky130_fd_sc_hd__o21a_1
X_4887_ _4910_/S vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__clkbuf_2
X_3907_ _6657_/Q _4262_/A _4264_/A _6656_/Q vssd1 vssd1 vccd1 vccd1 _3908_/D sky130_fd_sc_hd__a22o_1
X_6626_ _6799_/CLK _6626_/D vssd1 vssd1 vccd1 vccd1 _6626_/Q sky130_fd_sc_hd__dfxtp_1
X_3838_ _3850_/A _3849_/A _5214_/A _5214_/B vssd1 vssd1 vccd1 vccd1 _3839_/B sky130_fd_sc_hd__nand4_1
X_6557_ _6558_/CLK _6557_/D vssd1 vssd1 vccd1 vccd1 _6895_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3769_ _3769_/A _3769_/B _3769_/C vssd1 vssd1 vccd1 vccd1 _3769_/X sky130_fd_sc_hd__or3_1
XFILLER_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5508_ _6446_/Q _5652_/B vssd1 vssd1 vccd1 vccd1 _5508_/X sky130_fd_sc_hd__and2_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6488_ _6795_/CLK _6488_/D vssd1 vssd1 vccd1 vccd1 _6488_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5439_ _5439_/A _5439_/B vssd1 vssd1 vccd1 vccd1 _5440_/A sky130_fd_sc_hd__and2_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6551_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _6421_/Q _4812_/B vssd1 vssd1 vccd1 vccd1 _4811_/A sky130_fd_sc_hd__and2_1
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5790_ _6704_/Q _5755_/X _5789_/X _5773_/X vssd1 vssd1 vccd1 vccd1 _6704_/D sky130_fd_sc_hd__o211a_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4741_/A vssd1 vssd1 vccd1 vccd1 _6438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4672_ _4672_/A vssd1 vssd1 vccd1 vccd1 _6407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3623_ _3671_/A _3671_/B _3671_/C vssd1 vssd1 vccd1 vccd1 _3625_/B sky130_fd_sc_hd__nor3_1
X_6411_ _6789_/CLK _6411_/D vssd1 vssd1 vccd1 vccd1 _6411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6342_ _6789_/CLK _6342_/D vssd1 vssd1 vccd1 vccd1 _6342_/Q sky130_fd_sc_hd__dfxtp_1
X_3554_ _6651_/Q vssd1 vssd1 vccd1 vccd1 _3690_/B sky130_fd_sc_hd__clkbuf_2
X_3485_ _3485_/A vssd1 vssd1 vccd1 vccd1 _6320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6273_ _6273_/A _6283_/B vssd1 vssd1 vccd1 vccd1 _6273_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5224_ _5224_/A _5224_/B _5224_/C _5224_/D vssd1 vssd1 vccd1 vccd1 _5236_/A sky130_fd_sc_hd__or4_4
X_5155_ _5186_/A vssd1 vssd1 vccd1 vccd1 _5180_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5086_ _5086_/A vssd1 vssd1 vccd1 vccd1 _5109_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4106_ _4106_/A _4106_/B _4106_/C vssd1 vssd1 vccd1 vccd1 _4106_/Y sky130_fd_sc_hd__nand3_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4037_ _6663_/Q vssd1 vssd1 vccd1 vccd1 _4153_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _5969_/X _5985_/X _5987_/X vssd1 vssd1 vccd1 vccd1 _5988_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4939_ _6537_/Q _4939_/B vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__nor2_8
XFILLER_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6609_ _6667_/CLK _6609_/D vssd1 vssd1 vccd1 vccd1 _6609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3270_ _3274_/A vssd1 vssd1 vccd1 vccd1 _3270_/Y sky130_fd_sc_hd__inv_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6960_ _6960_/A _3261_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5911_ _6725_/Q _5888_/X _5910_/X _5904_/X vssd1 vssd1 vccd1 vccd1 _6725_/D sky130_fd_sc_hd__o211a_1
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5842_ _5619_/X _5841_/X _5842_/S vssd1 vssd1 vccd1 vccd1 _5842_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5773_ _5838_/A vssd1 vssd1 vccd1 vccd1 _5773_/X sky130_fd_sc_hd__clkbuf_2
X_4724_ _4735_/A vssd1 vssd1 vccd1 vccd1 _4733_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4655_ _6336_/Q _4655_/B vssd1 vssd1 vccd1 vccd1 _4656_/A sky130_fd_sc_hd__and2_1
Xinput60 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 _4928_/B sky130_fd_sc_hd__clkbuf_2
X_4586_ _4584_/Y _4555_/B _4585_/X vssd1 vssd1 vccd1 vccd1 _4607_/B sky130_fd_sc_hd__a21bo_1
X_3606_ _6654_/Q vssd1 vssd1 vccd1 vccd1 _3789_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6325_ _6554_/CLK _6325_/D vssd1 vssd1 vccd1 vccd1 _6325_/Q sky130_fd_sc_hd__dfxtp_1
X_3537_ _3534_/Y _3549_/B _3536_/X vssd1 vssd1 vccd1 vccd1 _3538_/B sky130_fd_sc_hd__o21ai_1
XFILLER_115_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3468_ _3468_/A vssd1 vssd1 vccd1 vccd1 _6312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6256_ _6806_/Q _6247_/X _6254_/Y _6255_/X vssd1 vssd1 vccd1 vccd1 _6806_/D sky130_fd_sc_hd__o211a_1
X_3399_ _3399_/A vssd1 vssd1 vccd1 vccd1 _6294_/D sky130_fd_sc_hd__clkbuf_1
X_5207_ _5243_/A _5207_/B _5207_/C vssd1 vssd1 vccd1 vccd1 _5208_/A sky130_fd_sc_hd__and3_1
X_6187_ _6785_/Q _5342_/X _6186_/X _6178_/X vssd1 vssd1 vccd1 vccd1 _6785_/D sky130_fd_sc_hd__o211a_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5138_ _5169_/A vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5069_ _6900_/A _5041_/X _5067_/X _5068_/X vssd1 vssd1 vccd1 vccd1 _6562_/D sky130_fd_sc_hd__o211a_1
XFILLER_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4440_ _4517_/A _4550_/C _6378_/Q _4368_/B vssd1 vssd1 vccd1 vccd1 _4442_/A sky130_fd_sc_hd__a22oi_1
XFILLER_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4371_ _4368_/X _4371_/B _6666_/Q _4371_/D vssd1 vssd1 vccd1 vccd1 _4371_/X sky130_fd_sc_hd__and4b_1
X_6110_ _6110_/A _6110_/B vssd1 vssd1 vccd1 vccd1 _6111_/A sky130_fd_sc_hd__and2_1
X_3322_ _6545_/Q _6544_/Q _6546_/Q vssd1 vssd1 vccd1 vccd1 _3323_/B sky130_fd_sc_hd__o21a_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3253_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3253_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6041_ _6490_/Q _6023_/X _6249_/A _6031_/X vssd1 vssd1 vccd1 vccd1 _6041_/X sky130_fd_sc_hd__a31o_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _3187_/A vssd1 vssd1 vccd1 vccd1 _3184_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6943_ _6943_/A _3240_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_81_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5825_ _5946_/A vssd1 vssd1 vccd1 vccd1 _5825_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5756_ _6700_/Q _5643_/X _5770_/S vssd1 vssd1 vccd1 vccd1 _5756_/X sky130_fd_sc_hd__mux2_1
X_4707_ _6367_/Q _4711_/B vssd1 vssd1 vccd1 vccd1 _4708_/A sky130_fd_sc_hd__and2_1
X_5687_ _5843_/A vssd1 vssd1 vccd1 vccd1 _5687_/X sky130_fd_sc_hd__buf_2
XFILLER_118_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4638_ _4638_/A _4642_/B vssd1 vssd1 vccd1 vccd1 _4638_/X sky130_fd_sc_hd__and2_1
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4569_ _4615_/B _4568_/X _3781_/X vssd1 vssd1 vccd1 vccd1 _4569_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6308_ _6522_/CLK _6308_/D vssd1 vssd1 vccd1 vccd1 _6308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6239_ _6802_/Q _6226_/X _6238_/Y _6235_/X vssd1 vssd1 vccd1 vccd1 _6802_/D sky130_fd_sc_hd__o211a_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3940_ _3940_/A _3940_/B vssd1 vssd1 vccd1 vccd1 _3959_/A sky130_fd_sc_hd__xnor2_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3871_ _5217_/A _6275_/A vssd1 vssd1 vccd1 vccd1 _3872_/A sky130_fd_sc_hd__and2_1
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6590_ _6667_/CLK _6590_/D vssd1 vssd1 vccd1 vccd1 _6590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5610_ _6471_/Q vssd1 vssd1 vccd1 vccd1 _5610_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5541_ _6673_/Q _5523_/X _5532_/X _5539_/X _5540_/X vssd1 vssd1 vccd1 vccd1 _6673_/D
+ sky130_fd_sc_hd__o221a_1
X_5472_ _5472_/A vssd1 vssd1 vccd1 vccd1 _6663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4423_ _4382_/A _4385_/B _4463_/A _4421_/X vssd1 vssd1 vccd1 vccd1 _4463_/B sky130_fd_sc_hd__o211ai_2
X_4354_ _4499_/A _4354_/B _4354_/C vssd1 vssd1 vccd1 vccd1 _4354_/X sky130_fd_sc_hd__and3_1
X_3305_ _3305_/A vssd1 vssd1 vccd1 vccd1 _3310_/A sky130_fd_sc_hd__buf_12
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4285_ _6665_/Q vssd1 vssd1 vccd1 vccd1 _4451_/A sky130_fd_sc_hd__clkbuf_2
X_6024_ _6487_/Q _6023_/X _6013_/X _6003_/X vssd1 vssd1 vccd1 vccd1 _6024_/X sky130_fd_sc_hd__a31o_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3237_/A vssd1 vssd1 vccd1 vccd1 _3236_/Y sky130_fd_sc_hd__inv_2
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6824__84 vssd1 vssd1 vccd1 vccd1 _6824__84/HI _6933_/A sky130_fd_sc_hd__conb_1
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6926_ _6926_/A _3218_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5808_ _5836_/A vssd1 vssd1 vccd1 vccd1 _5808_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6788_ _6809_/CLK _6788_/D vssd1 vssd1 vccd1 vccd1 _6788_/Q sky130_fd_sc_hd__dfxtp_1
X_5739_ _5838_/A vssd1 vssd1 vccd1 vccd1 _5739_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _4070_/A _4069_/X vssd1 vssd1 vccd1 vccd1 _4072_/A sky130_fd_sc_hd__or2b_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4972_ _6541_/Q _4972_/B vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__and2_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3923_ _4153_/C vssd1 vssd1 vccd1 vccd1 _4266_/A sky130_fd_sc_hd__buf_2
X_6711_ _6532_/Q _6711_/D vssd1 vssd1 vccd1 vccd1 _6711_/Q sky130_fd_sc_hd__dfxtp_1
X_6642_ _6667_/CLK _6642_/D vssd1 vssd1 vccd1 vccd1 _6642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3854_ _3854_/A vssd1 vssd1 vccd1 vccd1 _3855_/C sky130_fd_sc_hd__inv_2
XFILLER_32_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6573_ _6580_/CLK _6573_/D vssd1 vssd1 vccd1 vccd1 _6911_/A sky130_fd_sc_hd__dfxtp_1
X_3785_ _3785_/A vssd1 vssd1 vccd1 vccd1 _3786_/A sky130_fd_sc_hd__inv_2
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5524_ _6463_/Q vssd1 vssd1 vccd1 vccd1 _5524_/X sky130_fd_sc_hd__clkbuf_4
X_5455_ _6307_/Q _4149_/B _5466_/S vssd1 vssd1 vccd1 vccd1 _5456_/B sky130_fd_sc_hd__mux2_1
X_4406_ _6380_/Q vssd1 vssd1 vccd1 vccd1 _4579_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5386_ _5719_/A vssd1 vssd1 vccd1 vccd1 _5770_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_113_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ _4368_/A _4368_/B _6374_/Q _4433_/D vssd1 vssd1 vccd1 vccd1 _4337_/X sky130_fd_sc_hd__and4_1
X_6860__120 vssd1 vssd1 vccd1 vccd1 _6860__120/HI _6969_/A sky130_fd_sc_hd__conb_1
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4268_ _4268_/A _4270_/B vssd1 vssd1 vccd1 vccd1 _4269_/A sky130_fd_sc_hd__and2_1
XFILLER_101_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3219_ _3219_/A vssd1 vssd1 vccd1 vccd1 _3224_/A sky130_fd_sc_hd__buf_12
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6007_ _6742_/Q _5581_/X _6017_/S vssd1 vssd1 vccd1 vccd1 _6007_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4199_ _4227_/A _4270_/A _4058_/B _4228_/A vssd1 vssd1 vccd1 vccd1 _4201_/A sky130_fd_sc_hd__a22o_1
XFILLER_82_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6909_ _6909_/A _3199_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__ebufn_8
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3570_ _3659_/A _5214_/D _3551_/A _3569_/X vssd1 vssd1 vccd1 vccd1 _3591_/A sky130_fd_sc_hd__a31o_1
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5240_ _5240_/A vssd1 vssd1 vccd1 vccd1 _6587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6844__104 vssd1 vssd1 vccd1 vccd1 _6844__104/HI _6953_/A sky130_fd_sc_hd__conb_1
X_5171_ _5150_/X _5170_/X _5145_/X vssd1 vssd1 vccd1 vccd1 _5172_/C sky130_fd_sc_hd__a21o_1
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4122_ _4122_/A _4122_/B vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__or2_1
X_4053_ _4074_/A _4074_/B _4074_/C vssd1 vssd1 vccd1 vccd1 _4062_/B sky130_fd_sc_hd__nand3_1
XFILLER_110_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput3 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4955_ _5113_/A vssd1 vssd1 vccd1 vccd1 _5043_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3906_ _3998_/C vssd1 vssd1 vccd1 vccd1 _4264_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4886_ _6509_/Q _4880_/X _4881_/X input67/X vssd1 vssd1 vccd1 vccd1 _6509_/D sky130_fd_sc_hd__a22o_1
X_6625_ _6799_/CLK _6625_/D vssd1 vssd1 vccd1 vccd1 _6625_/Q sky130_fd_sc_hd__dfxtp_1
X_3837_ _3849_/A _3810_/B _3808_/C _3850_/A vssd1 vssd1 vccd1 vccd1 _3839_/A sky130_fd_sc_hd__a22o_1
X_3768_ _3769_/A _3769_/B _3769_/C vssd1 vssd1 vccd1 vccd1 _3785_/A sky130_fd_sc_hd__o21ai_2
X_6556_ _6558_/CLK _6556_/D vssd1 vssd1 vccd1 vccd1 _6894_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5507_ _5668_/B vssd1 vssd1 vccd1 vccd1 _5652_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6487_ _6795_/CLK _6487_/D vssd1 vssd1 vccd1 vccd1 _6487_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3699_ _3653_/B _3698_/Y _3596_/A _3755_/C vssd1 vssd1 vccd1 vccd1 _3741_/A sky130_fd_sc_hd__o211a_1
XFILLER_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5438_ _3879_/A _3849_/A _5448_/S vssd1 vssd1 vccd1 vccd1 _5439_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5369_ _5369_/A vssd1 vssd1 vccd1 vccd1 _6631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _6390_/Q _4744_/B vssd1 vssd1 vccd1 vccd1 _4741_/A sky130_fd_sc_hd__and2_1
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4671_ _6343_/Q _4677_/B vssd1 vssd1 vccd1 vccd1 _4672_/A sky130_fd_sc_hd__and2_1
X_6410_ _6789_/CLK _6410_/D vssd1 vssd1 vccd1 vccd1 _6410_/Q sky130_fd_sc_hd__dfxtp_1
X_3622_ _3622_/A _3622_/B _3622_/C vssd1 vssd1 vccd1 vccd1 _3671_/C sky130_fd_sc_hd__and3_1
X_6341_ _6789_/CLK _6341_/D vssd1 vssd1 vccd1 vccd1 _6341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3553_ _6652_/Q vssd1 vssd1 vccd1 vccd1 _3753_/A sky130_fd_sc_hd__clkbuf_2
X_3484_ _6320_/Q _6524_/Q _3484_/S vssd1 vssd1 vccd1 vccd1 _3485_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6272_ _6810_/Q _6267_/X _6271_/Y _6255_/X vssd1 vssd1 vccd1 vccd1 _6810_/D sky130_fd_sc_hd__o211a_1
XFILLER_115_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5223_ _5223_/A _5223_/B _5223_/C vssd1 vssd1 vccd1 vccd1 _5224_/D sky130_fd_sc_hd__or3_2
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5154_ _5154_/A vssd1 vssd1 vccd1 vccd1 _6576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4105_ _4106_/B _4106_/C _4106_/A vssd1 vssd1 vccd1 vccd1 _4105_/X sky130_fd_sc_hd__a21o_1
X_5085_ _5108_/A _5085_/B vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__or2_1
XFILLER_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4036_ _4036_/A _4057_/B _4036_/C vssd1 vssd1 vccd1 vccd1 _4074_/A sky130_fd_sc_hd__and3_1
XFILLER_25_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ _6480_/Q _6056_/B _5986_/X _5976_/X vssd1 vssd1 vccd1 vccd1 _5987_/X sky130_fd_sc_hd__a31o_1
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4938_ _6534_/Q _6533_/Q _6535_/Q vssd1 vssd1 vccd1 vccd1 _4939_/B sky130_fd_sc_hd__o21a_1
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4869_ _4929_/S vssd1 vssd1 vccd1 vccd1 _4870_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_30 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6608_ _6667_/CLK _6608_/D vssd1 vssd1 vccd1 vccd1 _6608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6539_ _6546_/CLK _6539_/D vssd1 vssd1 vccd1 vccd1 _6539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5910_ _5906_/X _5907_/X _5909_/X _5767_/X vssd1 vssd1 vccd1 vccd1 _5910_/X sky130_fd_sc_hd__a211o_1
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5841_ _6714_/Q _5621_/X _5841_/S vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__mux2_1
X_5772_ _6493_/Q _5734_/A _5699_/X _5771_/X _5743_/X vssd1 vssd1 vccd1 vccd1 _5772_/X
+ sky130_fd_sc_hd__a221o_1
X_4723_ _4723_/A vssd1 vssd1 vccd1 vccd1 _6430_/D sky130_fd_sc_hd__clkbuf_1
X_4654_ _4654_/A vssd1 vssd1 vccd1 vccd1 _6399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4585_ _4585_/A _4554_/A vssd1 vssd1 vccd1 vccd1 _4585_/X sky130_fd_sc_hd__or2b_1
Xinput50 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput61 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_4
X_3605_ _3650_/A _3605_/B _3605_/C _3660_/A vssd1 vssd1 vccd1 vccd1 _3660_/B sky130_fd_sc_hd__nand4_2
X_6324_ _6528_/CLK _6324_/D vssd1 vssd1 vccd1 vccd1 _6324_/Q sky130_fd_sc_hd__dfxtp_1
X_3536_ _6648_/Q _3762_/D _3534_/B _3661_/A vssd1 vssd1 vccd1 vccd1 _3536_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6255_ _6255_/A vssd1 vssd1 vccd1 vccd1 _6255_/X sky130_fd_sc_hd__buf_2
X_3467_ _6312_/Q _6516_/Q _3473_/S vssd1 vssd1 vccd1 vccd1 _3468_/A sky130_fd_sc_hd__mux2_1
X_5206_ _5181_/X _5205_/X _5088_/A vssd1 vssd1 vccd1 vccd1 _5207_/C sky130_fd_sc_hd__a21o_1
X_3398_ _3396_/X _3398_/B _3398_/C vssd1 vssd1 vccd1 vccd1 _3399_/A sky130_fd_sc_hd__and3b_1
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6186_ _6233_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _6186_/X sky130_fd_sc_hd__or2_1
XFILLER_96_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5137_ _6912_/A _5149_/B vssd1 vssd1 vccd1 vccd1 _5141_/B sky130_fd_sc_hd__or2_1
XFILLER_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5068_ _6136_/A vssd1 vssd1 vccd1 vccd1 _5068_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4019_ _4019_/A _4019_/B _4019_/C vssd1 vssd1 vccd1 vccd1 _4067_/C sky130_fd_sc_hd__and3_1
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4370_ _4368_/A _4433_/D _4393_/C _4479_/B vssd1 vssd1 vccd1 vccd1 _4371_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3321_ _5001_/A vssd1 vssd1 vccd1 vccd1 _6330_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3252_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6040_ _6040_/A vssd1 vssd1 vccd1 vccd1 _6249_/A sky130_fd_sc_hd__buf_2
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _3187_/A vssd1 vssd1 vccd1 vccd1 _3183_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6942_ _6942_/A _3239_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5824_ _5824_/A vssd1 vssd1 vccd1 vccd1 _5946_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5755_ _5797_/A vssd1 vssd1 vccd1 vccd1 _5755_/X sky130_fd_sc_hd__buf_2
X_4706_ _4706_/A vssd1 vssd1 vccd1 vccd1 _6422_/D sky130_fd_sc_hd__clkbuf_1
X_5686_ _5506_/X _5682_/X _5721_/S vssd1 vssd1 vccd1 vccd1 _5686_/X sky130_fd_sc_hd__mux2_1
X_4637_ _4637_/A _4637_/B _4637_/C vssd1 vssd1 vccd1 vccd1 _4640_/A sky130_fd_sc_hd__and3_1
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4568_ _4615_/A _4615_/C _4567_/Y vssd1 vssd1 vccd1 vccd1 _4568_/X sky130_fd_sc_hd__o21a_1
XFILLER_103_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4499_ _4499_/A _4636_/B _4499_/C vssd1 vssd1 vccd1 vccd1 _4499_/X sky130_fd_sc_hd__and3_1
X_6307_ _6522_/CLK _6307_/D vssd1 vssd1 vccd1 vccd1 _6307_/Q sky130_fd_sc_hd__dfxtp_1
X_3519_ _3729_/A vssd1 vssd1 vccd1 vccd1 _3552_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6238_ _6227_/X _6237_/Y _6230_/X vssd1 vssd1 vccd1 vccd1 _6238_/Y sky130_fd_sc_hd__o21ai_1
X_6169_ _6169_/A vssd1 vssd1 vccd1 vccd1 _6169_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3870_ _3870_/A vssd1 vssd1 vccd1 vccd1 _6352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5540_ _5707_/A vssd1 vssd1 vccd1 vccd1 _5540_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5471_ _5474_/A _5471_/B vssd1 vssd1 vccd1 vccd1 _5472_/A sky130_fd_sc_hd__and2_1
X_4422_ _4463_/A _4421_/X _4382_/A _4385_/B vssd1 vssd1 vccd1 vccd1 _4424_/B sky130_fd_sc_hd__a211o_1
XFILLER_113_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4353_ _4350_/A _4349_/B _4350_/Y _4352_/X vssd1 vssd1 vccd1 vccd1 _6386_/D sky130_fd_sc_hd__o211a_1
X_3304_ _3304_/A vssd1 vssd1 vccd1 vccd1 _3304_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4284_ _4284_/A vssd1 vssd1 vccd1 vccd1 _6382_/D sky130_fd_sc_hd__clkbuf_1
X_3235_ _3237_/A vssd1 vssd1 vccd1 vccd1 _3235_/Y sky130_fd_sc_hd__inv_2
X_6023_ _6023_/A vssd1 vssd1 vccd1 vccd1 _6023_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6925_ _6925_/A _3312_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6787_ _6809_/CLK _6787_/D vssd1 vssd1 vccd1 vccd1 _6787_/Q sky130_fd_sc_hd__dfxtp_1
X_3999_ _4123_/A _4116_/B _4000_/C _4057_/A vssd1 vssd1 vccd1 vccd1 _4036_/A sky130_fd_sc_hd__a22o_1
X_5807_ _5560_/X _5806_/X _5814_/S vssd1 vssd1 vccd1 vccd1 _5807_/X sky130_fd_sc_hd__mux2_1
X_5738_ _6260_/A _5734_/X _5735_/X _5737_/X _5695_/X vssd1 vssd1 vccd1 vccd1 _5738_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _6687_/Q _5668_/X _5669_/S vssd1 vssd1 vccd1 vccd1 _5670_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4971_ _4972_/B _4971_/B vssd1 vssd1 vccd1 vccd1 _6540_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3922_ _6353_/Q vssd1 vssd1 vccd1 vccd1 _4153_/C sky130_fd_sc_hd__clkbuf_2
X_6710_ _6809_/CLK _6710_/D vssd1 vssd1 vccd1 vccd1 _6710_/Q sky130_fd_sc_hd__dfxtp_1
X_6641_ _6667_/CLK _6641_/D vssd1 vssd1 vccd1 vccd1 _6641_/Q sky130_fd_sc_hd__dfxtp_1
X_3853_ _3853_/A _3853_/B vssd1 vssd1 vccd1 vccd1 _3854_/A sky130_fd_sc_hd__xnor2_1
XFILLER_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6572_ _6580_/CLK _6572_/D vssd1 vssd1 vccd1 vccd1 _6910_/A sky130_fd_sc_hd__dfxtp_1
X_3784_ _3828_/B _3780_/X _3826_/B vssd1 vssd1 vccd1 vccd1 _3804_/A sky130_fd_sc_hd__o21bai_1
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5523_ _6011_/A vssd1 vssd1 vccd1 vccd1 _5523_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5454_ _5454_/A vssd1 vssd1 vccd1 vccd1 _6658_/D sky130_fd_sc_hd__clkbuf_1
X_4405_ _4404_/B _4404_/C _4404_/A vssd1 vssd1 vccd1 vccd1 _4428_/C sky130_fd_sc_hd__a21o_1
X_5385_ _6637_/Q _6636_/Q _5778_/B vssd1 vssd1 vccd1 vccd1 _5719_/A sky130_fd_sc_hd__and3b_1
X_4336_ _6375_/Q vssd1 vssd1 vccd1 vccd1 _4433_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4267_ _4267_/A vssd1 vssd1 vccd1 vccd1 _6377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6006_ _6741_/Q _5984_/X _6005_/X _5999_/X vssd1 vssd1 vccd1 vccd1 _6741_/D sky130_fd_sc_hd__o211a_1
XFILLER_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3218_ _3218_/A vssd1 vssd1 vccd1 vccd1 _3218_/Y sky130_fd_sc_hd__inv_2
X_4198_ _4198_/A _4198_/B vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__or2_1
XFILLER_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ _6908_/A _3198_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__ebufn_8
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6883__143 vssd1 vssd1 vccd1 vccd1 _6883__143/HI _6992_/A sky130_fd_sc_hd__conb_1
XFILLER_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5170_ _6696_/Q _6728_/Q _6760_/Q _6792_/Q _5157_/X _5169_/X vssd1 vssd1 vccd1 vccd1
+ _5170_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4121_ _4121_/A _4121_/B _6355_/Q _6356_/Q vssd1 vssd1 vccd1 vccd1 _4122_/B sky130_fd_sc_hd__and4_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4052_ _4052_/A _4052_/B _4052_/C vssd1 vssd1 vccd1 vccd1 _4074_/C sky130_fd_sc_hd__nand3_1
Xinput4 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4954_ _6535_/Q vssd1 vssd1 vccd1 vccd1 _5113_/A sky130_fd_sc_hd__buf_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3905_ _4083_/A vssd1 vssd1 vccd1 vccd1 _3941_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4885_ _6508_/Q _4880_/X _4881_/X input66/X vssd1 vssd1 vccd1 vccd1 _6508_/D sky130_fd_sc_hd__a22o_1
X_6624_ _6799_/CLK _6624_/D vssd1 vssd1 vccd1 vccd1 _6624_/Q sky130_fd_sc_hd__dfxtp_1
X_3836_ _3836_/A vssd1 vssd1 vccd1 vccd1 _3850_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3767_ _3797_/A _3767_/B vssd1 vssd1 vccd1 vccd1 _3769_/C sky130_fd_sc_hd__xnor2_1
XFILLER_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6555_ _6558_/CLK _6555_/D vssd1 vssd1 vccd1 vccd1 _6893_/A sky130_fd_sc_hd__dfxtp_1
X_5506_ _6462_/Q vssd1 vssd1 vccd1 vccd1 _5506_/X sky130_fd_sc_hd__buf_2
X_6486_ _6763_/CLK _6486_/D vssd1 vssd1 vccd1 vccd1 _6486_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3698_ _3698_/A _3698_/B vssd1 vssd1 vccd1 vccd1 _3698_/Y sky130_fd_sc_hd__nor2_1
X_5437_ _5437_/A vssd1 vssd1 vccd1 vccd1 _6653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5368_ _6631_/Q _5372_/B vssd1 vssd1 vccd1 vccd1 _5369_/A sky130_fd_sc_hd__and2_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5299_ _6613_/Q _5305_/B vssd1 vssd1 vccd1 vccd1 _5300_/A sky130_fd_sc_hd__and2_1
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4319_ _4319_/A _4319_/B vssd1 vssd1 vccd1 vccd1 _4320_/B sky130_fd_sc_hd__and2_1
XFILLER_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6867__127 vssd1 vssd1 vccd1 vccd1 _6867__127/HI _6976_/A sky130_fd_sc_hd__conb_1
XFILLER_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _4670_/A vssd1 vssd1 vccd1 vccd1 _6406_/D sky130_fd_sc_hd__clkbuf_1
X_3621_ _3622_/B _3622_/C _3622_/A vssd1 vssd1 vccd1 vccd1 _3671_/B sky130_fd_sc_hd__a21oi_1
X_3552_ _3552_/A _5217_/B vssd1 vssd1 vccd1 vccd1 _3559_/A sky130_fd_sc_hd__nand2_1
X_6340_ _6789_/CLK _6340_/D vssd1 vssd1 vccd1 vccd1 _6340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6271_ _6268_/X _6270_/Y _6264_/X vssd1 vssd1 vccd1 vccd1 _6271_/Y sky130_fd_sc_hd__o21ai_1
X_3483_ _3483_/A vssd1 vssd1 vccd1 vccd1 _6319_/D sky130_fd_sc_hd__clkbuf_1
X_5222_ _6315_/Q _6314_/Q _6313_/Q _6312_/Q vssd1 vssd1 vccd1 vccd1 _5223_/C sky130_fd_sc_hd__or4_1
X_5153_ _5160_/A _5153_/B _5153_/C vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__and3_1
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4104_ _3889_/A _4275_/A _4060_/B _4103_/X vssd1 vssd1 vccd1 vccd1 _4106_/A sky130_fd_sc_hd__a31o_1
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5084_ _6682_/Q _6714_/Q _6746_/Q _6778_/Q _5083_/X _5063_/X vssd1 vssd1 vccd1 vccd1
+ _5085_/B sky130_fd_sc_hd__mux4_1
XFILLER_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4035_ _4067_/C vssd1 vssd1 vccd1 vccd1 _4035_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _6040_/A vssd1 vssd1 vccd1 vccd1 _5986_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ _4935_/X _4936_/X _6543_/Q vssd1 vssd1 vccd1 vccd1 _5017_/B sky130_fd_sc_hd__a21o_1
X_4868_ _3362_/Y _4867_/B _4867_/Y _3361_/X _3632_/A vssd1 vssd1 vccd1 vccd1 _4929_/S
+ sky130_fd_sc_hd__a2111o_4
XANTENNA_31 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_20 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6607_ _6667_/CLK _6607_/D vssd1 vssd1 vccd1 vccd1 _6607_/Q sky130_fd_sc_hd__dfxtp_1
X_3819_ _3819_/A _3855_/A vssd1 vssd1 vccd1 vccd1 _3833_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4799_ _4799_/A vssd1 vssd1 vccd1 vccd1 _6464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6538_ _6546_/CLK _6538_/D vssd1 vssd1 vccd1 vccd1 _6538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6469_ _6763_/CLK _6469_/D vssd1 vssd1 vccd1 vccd1 _6469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5840_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5840_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5771_ _6477_/Q _5770_/X _5771_/S vssd1 vssd1 vccd1 vccd1 _5771_/X sky130_fd_sc_hd__mux2_1
X_4722_ _6382_/Q _4722_/B vssd1 vssd1 vccd1 vccd1 _4723_/A sky130_fd_sc_hd__and2_1
Xinput40 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_2
X_4653_ _6335_/Q _4655_/B vssd1 vssd1 vccd1 vccd1 _4654_/A sky130_fd_sc_hd__and2_1
X_4584_ _4584_/A vssd1 vssd1 vccd1 vccd1 _4584_/Y sky130_fd_sc_hd__inv_2
Xinput51 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_4
X_3604_ _6300_/Q vssd1 vssd1 vccd1 vccd1 _3605_/B sky130_fd_sc_hd__clkbuf_2
Xinput62 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6323_ _6528_/CLK _6323_/D vssd1 vssd1 vccd1 vccd1 _6323_/Q sky130_fd_sc_hd__dfxtp_1
X_3535_ _3661_/A _3762_/D vssd1 vssd1 vccd1 vccd1 _3549_/B sky130_fd_sc_hd__nand2_1
X_3466_ _3466_/A vssd1 vssd1 vccd1 vccd1 _6311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6254_ _6248_/X _6253_/Y _6244_/X vssd1 vssd1 vccd1 vccd1 _6254_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_107_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5205_ _6702_/Q _6734_/Q _6766_/Q _6798_/Q _5188_/X _5014_/X vssd1 vssd1 vccd1 vccd1
+ _5205_/X sky130_fd_sc_hd__mux4_1
X_3397_ _6293_/Q _3396_/C _6294_/Q vssd1 vssd1 vccd1 vccd1 _3398_/C sky130_fd_sc_hd__a21o_1
X_6185_ _6784_/Q _5342_/X _6184_/X _6178_/X vssd1 vssd1 vccd1 vccd1 _6784_/D sky130_fd_sc_hd__o211a_1
X_5136_ _5136_/A vssd1 vssd1 vccd1 vccd1 _6573_/D sky130_fd_sc_hd__clkbuf_1
X_5067_ _5047_/X _5065_/X _5066_/X _5055_/X vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__a31o_1
X_4018_ _4019_/B _4019_/C _4019_/A vssd1 vssd1 vccd1 vccd1 _4067_/B sky130_fd_sc_hd__a21oi_1
XFILLER_53_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5969_ _6029_/A vssd1 vssd1 vccd1 vccd1 _5969_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3320_ _3632_/A vssd1 vssd1 vccd1 vccd1 _5001_/A sky130_fd_sc_hd__buf_4
XFILLER_98_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3251_/Y sky130_fd_sc_hd__inv_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3182_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3187_/A sky130_fd_sc_hd__buf_2
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6941_ _6941_/A _3237_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5823_ _6710_/Q _5797_/X _5822_/X _5810_/X vssd1 vssd1 vccd1 vccd1 _6710_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5754_ _6699_/Q _5718_/X _5753_/X _5739_/X vssd1 vssd1 vccd1 vccd1 _6699_/D sky130_fd_sc_hd__o211a_1
X_4705_ _6366_/Q _4711_/B vssd1 vssd1 vccd1 vccd1 _4706_/A sky130_fd_sc_hd__and2_1
X_5685_ _5771_/S vssd1 vssd1 vccd1 vccd1 _5721_/S sky130_fd_sc_hd__clkbuf_2
X_4636_ _4636_/A _4636_/B vssd1 vssd1 vccd1 vccd1 _4637_/C sky130_fd_sc_hd__nand2_1
X_4567_ _4566_/A _4566_/D _4566_/C vssd1 vssd1 vccd1 vccd1 _4567_/Y sky130_fd_sc_hd__o21bai_1
X_6306_ _6522_/CLK _6306_/D vssd1 vssd1 vccd1 vccd1 _6306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4498_ _4595_/D vssd1 vssd1 vccd1 vccd1 _4636_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3518_ _3650_/A vssd1 vssd1 vccd1 vccd1 _3729_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3449_ _6304_/Q _6508_/Q _3451_/S vssd1 vssd1 vccd1 vccd1 _3450_/A sky130_fd_sc_hd__mux2_1
X_6237_ _6237_/A _6243_/B vssd1 vssd1 vccd1 vccd1 _6237_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6777_/Q _6156_/X _6167_/X _6165_/X vssd1 vssd1 vccd1 vccd1 _6777_/D sky130_fd_sc_hd__o211a_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5119_ _5181_/A vssd1 vssd1 vccd1 vccd1 _5119_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6099_ _6110_/A _6099_/B vssd1 vssd1 vccd1 vccd1 _6100_/A sky130_fd_sc_hd__and2_1
XFILLER_72_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5470_ _6311_/Q _4242_/A _5483_/S vssd1 vssd1 vccd1 vccd1 _5471_/B sky130_fd_sc_hd__mux2_1
X_4421_ _4420_/A _4420_/B _4420_/C vssd1 vssd1 vccd1 vccd1 _4421_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4352_ _6136_/A vssd1 vssd1 vccd1 vccd1 _4352_/X sky130_fd_sc_hd__buf_6
XFILLER_113_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3303_ _3304_/A vssd1 vssd1 vccd1 vccd1 _3303_/Y sky130_fd_sc_hd__inv_2
X_4283_ _4283_/A _4300_/B _5008_/B vssd1 vssd1 vccd1 vccd1 _4284_/A sky130_fd_sc_hd__and3_1
X_3234_ _3237_/A vssd1 vssd1 vccd1 vccd1 _3234_/Y sky130_fd_sc_hd__inv_2
X_6022_ _6745_/Q _5610_/X _6044_/S vssd1 vssd1 vccd1 vccd1 _6022_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924_ _6924_/A _3217_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__ebufn_8
XFILLER_82_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6786_ _6789_/CLK _6786_/D vssd1 vssd1 vccd1 vccd1 _6786_/Q sky130_fd_sc_hd__dfxtp_1
X_3998_ _4147_/A _4085_/B _3998_/C _3998_/D vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__nand4_2
X_5806_ _6708_/Q _5561_/X _5813_/S vssd1 vssd1 vccd1 vccd1 _5806_/X sky130_fd_sc_hd__mux2_1
X_5737_ _5602_/X _5736_/X _5757_/S vssd1 vssd1 vccd1 vccd1 _5737_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5668_ _6461_/Q _5668_/B vssd1 vssd1 vccd1 vccd1 _5668_/X sky130_fd_sc_hd__and2_2
X_4619_ _4619_/A vssd1 vssd1 vccd1 vccd1 _6394_/D sky130_fd_sc_hd__clkbuf_1
X_5599_ _6257_/A _5589_/X _5578_/X _5567_/X vssd1 vssd1 vccd1 vccd1 _5599_/X sky130_fd_sc_hd__a31o_1
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4970_ _6540_/Q _4968_/A _4931_/X vssd1 vssd1 vccd1 vccd1 _4971_/B sky130_fd_sc_hd__o21ai_1
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3921_ _4013_/A _4264_/A vssd1 vssd1 vccd1 vccd1 _3921_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6640_ _6532_/Q _6640_/D vssd1 vssd1 vccd1 vccd1 _6640_/Q sky130_fd_sc_hd__dfxtp_1
X_3852_ _3840_/A _3839_/A _3839_/B _3851_/X vssd1 vssd1 vccd1 vccd1 _3853_/B sky130_fd_sc_hd__a31o_1
XFILLER_20_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6571_ _6586_/CLK _6571_/D vssd1 vssd1 vccd1 vccd1 _6909_/A sky130_fd_sc_hd__dfxtp_1
X_5522_ _6672_/Q _3357_/X _5521_/X _5100_/X vssd1 vssd1 vccd1 vccd1 _6672_/D sky130_fd_sc_hd__o211a_1
X_3783_ _3828_/B _3780_/X _3782_/Y vssd1 vssd1 vccd1 vccd1 _6344_/D sky130_fd_sc_hd__a21oi_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5453_ _5456_/A _5453_/B vssd1 vssd1 vccd1 vccd1 _5454_/A sky130_fd_sc_hd__and2_1
X_4404_ _4404_/A _4404_/B _4404_/C vssd1 vssd1 vccd1 vccd1 _4428_/B sky130_fd_sc_hd__nand3_4
X_5384_ _6640_/Q _6639_/Q _6638_/Q _5509_/D vssd1 vssd1 vccd1 vccd1 _5778_/B sky130_fd_sc_hd__nor4_2
XFILLER_113_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4335_ _6667_/Q vssd1 vssd1 vccd1 vccd1 _4368_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4266_ _4266_/A _4270_/B vssd1 vssd1 vccd1 vccd1 _4267_/A sky130_fd_sc_hd__and2_1
XFILLER_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3217_ _3218_/A vssd1 vssd1 vccd1 vccd1 _3217_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6005_ _6001_/X _6002_/X _6004_/X vssd1 vssd1 vccd1 vccd1 _6005_/X sky130_fd_sc_hd__a21o_1
X_4197_ _4195_/X _4196_/Y _6067_/A vssd1 vssd1 vccd1 vccd1 _6369_/D sky130_fd_sc_hd__a21oi_1
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6907_ _6907_/A _3197_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__ebufn_8
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6769_ _6789_/CLK _6769_/D vssd1 vssd1 vccd1 vccd1 _6769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4120_ _3944_/A _6355_/Q _6356_/Q _3944_/B vssd1 vssd1 vccd1 vccd1 _4122_/A sky130_fd_sc_hd__a22oi_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4051_ _4052_/B _4052_/C _4052_/A vssd1 vssd1 vccd1 vccd1 _4074_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput5 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4953_ _4953_/A vssd1 vssd1 vccd1 vccd1 _6534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3904_ _6658_/Q vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__clkbuf_2
X_6623_ _6799_/CLK _6623_/D vssd1 vssd1 vccd1 vccd1 _6623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4884_ _6507_/Q _4880_/X _4881_/X input65/X vssd1 vssd1 vccd1 vccd1 _6507_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3835_ _3835_/A vssd1 vssd1 vccd1 vccd1 _3849_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6554_ _6554_/CLK _6554_/D vssd1 vssd1 vccd1 vccd1 _6554_/Q sky130_fd_sc_hd__dfxtp_1
X_3766_ _3766_/A _3798_/A vssd1 vssd1 vccd1 vccd1 _3767_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6485_ _6763_/CLK _6485_/D vssd1 vssd1 vccd1 vccd1 _6485_/Q sky130_fd_sc_hd__dfxtp_4
X_5505_ _5620_/A vssd1 vssd1 vccd1 vccd1 _5505_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3697_ _3696_/A _3696_/B _3696_/C vssd1 vssd1 vccd1 vccd1 _3703_/C sky130_fd_sc_hd__a21o_1
X_5436_ _5439_/A _5436_/B vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__and2_1
X_5367_ _5971_/A _5364_/X _5331_/X vssd1 vssd1 vccd1 vccd1 _6630_/D sky130_fd_sc_hd__o21a_1
XFILLER_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5298_ _5298_/A vssd1 vssd1 vccd1 vccd1 _6612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4318_ _4319_/A _4319_/B vssd1 vssd1 vccd1 vccd1 _4320_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4249_ _4249_/A _4249_/B vssd1 vssd1 vccd1 vccd1 _4249_/X sky130_fd_sc_hd__or2_1
XFILLER_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6850__110 vssd1 vssd1 vccd1 vccd1 _6850__110/HI _6959_/A sky130_fd_sc_hd__conb_1
X_3620_ _3620_/A _3639_/C vssd1 vssd1 vccd1 vccd1 _3622_/A sky130_fd_sc_hd__xnor2_1
X_3551_ _3551_/A _3551_/B vssd1 vssd1 vccd1 vccd1 _3571_/A sky130_fd_sc_hd__xnor2_1
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6270_ _6270_/A _6283_/B vssd1 vssd1 vccd1 vccd1 _6270_/Y sky130_fd_sc_hd__nand2_1
X_3482_ _6319_/Q _6523_/Q _3484_/S vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5221_ _6327_/Q _6326_/Q _6325_/Q _6324_/Q vssd1 vssd1 vccd1 vccd1 _5223_/B sky130_fd_sc_hd__or4_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5152_ _5150_/X _5151_/X _5145_/X vssd1 vssd1 vccd1 vccd1 _5153_/C sky130_fd_sc_hd__a21o_1
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4103_ _4103_/A _4273_/A _4103_/C vssd1 vssd1 vccd1 vccd1 _4103_/X sky130_fd_sc_hd__and3_1
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5083_ _6533_/Q vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__buf_2
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4034_ _3889_/A _4273_/A _4017_/B _4033_/X vssd1 vssd1 vccd1 vccd1 _4065_/A sky130_fd_sc_hd__a31oi_2
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5985_ _6738_/Q _5542_/X _5990_/S vssd1 vssd1 vccd1 vccd1 _5985_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4936_ _6542_/Q _6541_/Q _6540_/Q vssd1 vssd1 vccd1 vccd1 _4936_/X sky130_fd_sc_hd__and3_1
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_21 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4867_ _6330_/Q _4867_/B vssd1 vssd1 vccd1 vccd1 _4867_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_10 _3325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6606_ _6667_/CLK _6606_/D vssd1 vssd1 vccd1 vccd1 _6606_/Q sky130_fd_sc_hd__dfxtp_1
X_3818_ _3818_/A _3818_/B vssd1 vssd1 vccd1 vccd1 _3855_/A sky130_fd_sc_hd__nor2_1
XFILLER_122_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6537_ _6586_/CLK _6537_/D vssd1 vssd1 vccd1 vccd1 _6537_/Q sky130_fd_sc_hd__dfxtp_2
X_4798_ _6416_/Q _4800_/B vssd1 vssd1 vccd1 vccd1 _4799_/A sky130_fd_sc_hd__and2_1
X_3749_ _3749_/A _3749_/B vssd1 vssd1 vccd1 vccd1 _6343_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6468_ _6763_/CLK _6468_/D vssd1 vssd1 vccd1 vccd1 _6468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6399_ _6789_/CLK _6399_/D vssd1 vssd1 vccd1 vccd1 _6399_/Q sky130_fd_sc_hd__dfxtp_1
X_5419_ _5422_/A _5419_/B vssd1 vssd1 vccd1 vccd1 _5420_/A sky130_fd_sc_hd__and2_1
XFILLER_121_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5770_ _6703_/Q _5668_/X _5770_/S vssd1 vssd1 vccd1 vccd1 _5770_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4721_/A vssd1 vssd1 vccd1 vccd1 _6429_/D sky130_fd_sc_hd__clkbuf_1
X_4652_ _4652_/A vssd1 vssd1 vccd1 vccd1 _6398_/D sky130_fd_sc_hd__clkbuf_1
X_3603_ _3650_/A _3789_/D _3605_/C _3660_/A vssd1 vssd1 vccd1 vccd1 _3641_/A sky130_fd_sc_hd__a22o_1
Xinput30 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _3325_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput52 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 _4906_/B sky130_fd_sc_hd__clkbuf_1
X_4583_ _4583_/A _4583_/B vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__xnor2_1
Xinput41 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_2
Xinput63 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_2
X_6322_ _6531_/CLK _6322_/D vssd1 vssd1 vccd1 vccd1 _6322_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6531_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_3534_ _3616_/A _3534_/B vssd1 vssd1 vccd1 vccd1 _3534_/Y sky130_fd_sc_hd__nand2_1
X_3465_ _6311_/Q _6515_/Q _3473_/S vssd1 vssd1 vccd1 vccd1 _3466_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6253_ _6253_/A _6263_/B vssd1 vssd1 vccd1 vccd1 _6253_/Y sky130_fd_sc_hd__nand2_1
X_5204_ _6923_/A _5209_/B vssd1 vssd1 vccd1 vccd1 _5207_/B sky130_fd_sc_hd__or2_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3396_ _6294_/Q _6293_/Q _3396_/C vssd1 vssd1 vccd1 vccd1 _3396_/X sky130_fd_sc_hd__and3_1
X_6184_ _6229_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _6184_/X sky130_fd_sc_hd__or2_1
XFILLER_123_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5135_ _5160_/A _5135_/B _5135_/C vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__and3_1
XFILLER_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5066_ _6807_/Q _5078_/B vssd1 vssd1 vccd1 vccd1 _5066_/X sky130_fd_sc_hd__or2_1
XFILLER_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4017_ _4017_/A _4017_/B vssd1 vssd1 vccd1 vccd1 _4019_/A sky130_fd_sc_hd__xnor2_1
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5968_ _6023_/A _6269_/A vssd1 vssd1 vccd1 vccd1 _6029_/A sky130_fd_sc_hd__nand2_2
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4919_ _4919_/A _4919_/B vssd1 vssd1 vccd1 vccd1 _4919_/X sky130_fd_sc_hd__and2_1
XFILLER_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5899_ _5871_/X _5897_/X _5898_/X _5767_/X vssd1 vssd1 vccd1 vccd1 _5899_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3250_/A vssd1 vssd1 vccd1 vccd1 _3255_/A sky130_fd_sc_hd__buf_12
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3305_/A vssd1 vssd1 vccd1 vccd1 _3313_/A sky130_fd_sc_hd__buf_12
XFILLER_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6940_ _6940_/A _3236_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_81_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5822_ _6484_/Q _5812_/X _5821_/X _5808_/X _5815_/X vssd1 vssd1 vccd1 vccd1 _5822_/X
+ sky130_fd_sc_hd__a221o_1
X_5753_ _6273_/A _5734_/X _5735_/X _5752_/X _5743_/X vssd1 vssd1 vccd1 vccd1 _5753_/X
+ sky130_fd_sc_hd__a221o_1
X_4704_ _4704_/A vssd1 vssd1 vccd1 vccd1 _6421_/D sky130_fd_sc_hd__clkbuf_1
X_5684_ _5700_/A _6059_/A vssd1 vssd1 vccd1 vccd1 _5771_/S sky130_fd_sc_hd__or2_2
X_4635_ _4630_/A _4634_/Y _4630_/B vssd1 vssd1 vccd1 vccd1 _4635_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4566_ _4566_/A _4566_/B _4566_/C _4566_/D vssd1 vssd1 vccd1 vccd1 _4615_/C sky130_fd_sc_hd__or4_1
X_3517_ _6650_/Q vssd1 vssd1 vccd1 vccd1 _3650_/A sky130_fd_sc_hd__clkbuf_2
X_6305_ _6504_/CLK _6305_/D vssd1 vssd1 vccd1 vccd1 _6305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4497_ _6380_/Q vssd1 vssd1 vccd1 vccd1 _4595_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6236_ _6801_/Q _6226_/X _6234_/Y _6235_/X vssd1 vssd1 vccd1 vccd1 _6801_/D sky130_fd_sc_hd__o211a_1
X_3448_ _3448_/A vssd1 vssd1 vccd1 vccd1 _6303_/D sky130_fd_sc_hd__clkbuf_1
X_3379_ _5193_/A vssd1 vssd1 vccd1 vccd1 _5412_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6263_/A _6167_/B vssd1 vssd1 vccd1 vccd1 _6167_/X sky130_fd_sc_hd__or2_1
X_5118_ _6909_/A _5118_/B vssd1 vssd1 vccd1 vccd1 _5122_/B sky130_fd_sc_hd__or2_1
XFILLER_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6098_ _6758_/Q _6080_/X _6097_/X _6076_/X vssd1 vssd1 vccd1 vccd1 _6099_/B sky130_fd_sc_hd__a22o_1
X_5049_ _6533_/Q vssd1 vssd1 vccd1 vccd1 _5049_/X sky130_fd_sc_hd__buf_2
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4420_ _4420_/A _4420_/B _4420_/C vssd1 vssd1 vccd1 vccd1 _4463_/A sky130_fd_sc_hd__nand3_2
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4351_ _5458_/A vssd1 vssd1 vccd1 vccd1 _6136_/A sky130_fd_sc_hd__clkbuf_8
X_3302_ _3304_/A vssd1 vssd1 vccd1 vccd1 _3302_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4282_ _4373_/D vssd1 vssd1 vccd1 vccd1 _4300_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6021_ _6048_/S vssd1 vssd1 vccd1 vccd1 _6044_/S sky130_fd_sc_hd__clkbuf_2
X_3233_ _3237_/A vssd1 vssd1 vccd1 vccd1 _3233_/Y sky130_fd_sc_hd__inv_2
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6923_ _6923_/A _3216_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__ebufn_8
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6785_ _6799_/CLK _6785_/D vssd1 vssd1 vccd1 vccd1 _6785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5805_ _6707_/Q _5797_/X _5804_/X _5773_/X vssd1 vssd1 vccd1 vccd1 _6707_/D sky130_fd_sc_hd__o211a_1
X_3997_ _4121_/A vssd1 vssd1 vccd1 vccd1 _4147_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5736_ _6696_/Q _5603_/X _5751_/S vssd1 vssd1 vccd1 vccd1 _5736_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5667_ _6477_/Q vssd1 vssd1 vccd1 vccd1 _5667_/X sky130_fd_sc_hd__clkbuf_2
X_4618_ _4616_/X _4618_/B vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__and2b_1
XFILLER_123_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5598_ _6485_/Q vssd1 vssd1 vccd1 vccd1 _6257_/A sky130_fd_sc_hd__clkbuf_4
X_4549_ _4622_/A _4371_/B _4512_/B _4576_/B vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__a22oi_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6219_ _6797_/Q _6207_/X _6218_/X _6216_/X vssd1 vssd1 vccd1 vccd1 _6797_/D sky130_fd_sc_hd__o211a_1
XFILLER_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3920_ _3957_/C _3920_/B vssd1 vssd1 vccd1 vccd1 _3927_/A sky130_fd_sc_hd__or2_1
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3851_ _3851_/A _3855_/B vssd1 vssd1 vccd1 vccd1 _3851_/X sky130_fd_sc_hd__and2_1
XFILLER_20_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6570_ _6570_/CLK _6570_/D vssd1 vssd1 vccd1 vccd1 _6908_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3782_ _3828_/B _3780_/X _3781_/X vssd1 vssd1 vccd1 vccd1 _3782_/Y sky130_fd_sc_hd__o21ai_1
X_5521_ _5505_/X _5515_/X _5520_/X vssd1 vssd1 vccd1 vccd1 _5521_/X sky130_fd_sc_hd__a21o_1
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5452_ _6306_/Q _3941_/A _5466_/S vssd1 vssd1 vccd1 vccd1 _5453_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5383_ _5383_/A _5668_/B vssd1 vssd1 vccd1 vccd1 _5509_/D sky130_fd_sc_hd__nand2_1
X_4403_ _4429_/A _4450_/B _4429_/C vssd1 vssd1 vccd1 vccd1 _4404_/C sky130_fd_sc_hd__a21o_1
X_4334_ _6668_/Q vssd1 vssd1 vccd1 vccd1 _4368_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4265_ _4265_/A vssd1 vssd1 vccd1 vccd1 _6376_/D sky130_fd_sc_hd__clkbuf_1
X_6004_ _6483_/Q _5996_/X _5986_/X _6003_/X vssd1 vssd1 vccd1 vccd1 _6004_/X sky130_fd_sc_hd__a31o_1
X_3216_ _3218_/A vssd1 vssd1 vccd1 vccd1 _3216_/Y sky130_fd_sc_hd__inv_2
X_4196_ _4218_/B _4195_/B _4220_/D vssd1 vssd1 vccd1 vccd1 _4196_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6906_ _6906_/A _3196_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__ebufn_8
XFILLER_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6768_ _6789_/CLK _6768_/D vssd1 vssd1 vccd1 vccd1 _6768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5719_ _5719_/A vssd1 vssd1 vccd1 vccd1 _5751_/S sky130_fd_sc_hd__buf_2
X_6699_ _6809_/CLK _6699_/D vssd1 vssd1 vccd1 vccd1 _6699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _4093_/A _4093_/B vssd1 vssd1 vccd1 vccd1 _4052_/A sky130_fd_sc_hd__xor2_1
XFILLER_83_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput6 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
XFILLER_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4952_ _4950_/X _5239_/B _4952_/C vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__and3b_1
X_3903_ _6657_/Q _6656_/Q _4039_/D _3998_/C vssd1 vssd1 vccd1 vccd1 _3928_/A sky130_fd_sc_hd__and4_1
X_4883_ _6506_/Q _4880_/X _4881_/X input64/X vssd1 vssd1 vccd1 vccd1 _6506_/D sky130_fd_sc_hd__a22o_1
X_6622_ _6799_/CLK _6622_/D vssd1 vssd1 vccd1 vccd1 _6622_/Q sky130_fd_sc_hd__dfxtp_1
X_3834_ _3811_/A _3811_/B _3809_/B vssd1 vssd1 vccd1 vccd1 _3840_/A sky130_fd_sc_hd__o21ai_2
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6553_ _6580_/CLK _6553_/D vssd1 vssd1 vccd1 vccd1 _6892_/A sky130_fd_sc_hd__dfxtp_1
X_3765_ _3765_/A _3765_/B vssd1 vssd1 vccd1 vccd1 _3798_/A sky130_fd_sc_hd__and2_1
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5504_ _5957_/C _6040_/A vssd1 vssd1 vccd1 vccd1 _5620_/A sky130_fd_sc_hd__nand2_2
X_6484_ _6763_/CLK _6484_/D vssd1 vssd1 vccd1 vccd1 _6484_/Q sky130_fd_sc_hd__dfxtp_4
X_3696_ _3696_/A _3696_/B _3696_/C vssd1 vssd1 vccd1 vccd1 _3703_/B sky130_fd_sc_hd__nand3_2
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5435_ _5214_/C _3810_/A _5448_/S vssd1 vssd1 vccd1 vccd1 _5436_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5366_ _6630_/Q vssd1 vssd1 vccd1 vccd1 _5971_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5297_ _6612_/Q _5305_/B vssd1 vssd1 vccd1 vccd1 _5298_/A sky130_fd_sc_hd__and2_1
X_4317_ _4354_/B _4315_/X _4316_/X vssd1 vssd1 vccd1 vccd1 _4319_/B sky130_fd_sc_hd__a21bo_1
XFILLER_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4248_ _4247_/A _4247_/B _4247_/C vssd1 vssd1 vccd1 vccd1 _4249_/B sky130_fd_sc_hd__a21oi_1
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4179_ _4227_/A _4116_/B _4180_/D _4228_/A vssd1 vssd1 vccd1 vccd1 _4181_/A sky130_fd_sc_hd__a22oi_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3550_ _3616_/A _3722_/B vssd1 vssd1 vccd1 vccd1 _3551_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220_ _6323_/Q _6322_/Q _6321_/Q _6320_/Q vssd1 vssd1 vccd1 vccd1 _5223_/A sky130_fd_sc_hd__or4_1
X_3481_ _3481_/A vssd1 vssd1 vccd1 vccd1 _6318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5151_ _6693_/Q _6725_/Q _6757_/Q _6789_/Q _5126_/X _5138_/X vssd1 vssd1 vccd1 vccd1
+ _5151_/X sky130_fd_sc_hd__mux4_2
XFILLER_123_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5082_ _5113_/A vssd1 vssd1 vccd1 vccd1 _5108_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_57_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4102_ _4230_/D vssd1 vssd1 vccd1 vccd1 _4275_/A sky130_fd_sc_hd__buf_2
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4033_ _4103_/A _4270_/A _4033_/C vssd1 vssd1 vccd1 vccd1 _4033_/X sky130_fd_sc_hd__and3_1
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ _6011_/A vssd1 vssd1 vccd1 vccd1 _5984_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4935_ _6539_/Q _6538_/Q vssd1 vssd1 vccd1 vccd1 _4935_/X sky130_fd_sc_hd__or2_1
X_4866_ _6332_/Q _6333_/Q vssd1 vssd1 vccd1 vccd1 _4867_/B sky130_fd_sc_hd__or2_2
XANTENNA_11 _3327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_22 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6605_ _6667_/CLK _6605_/D vssd1 vssd1 vccd1 vccd1 _6605_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_33 _3325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3817_ _3818_/A _3818_/B vssd1 vssd1 vccd1 vccd1 _3819_/A sky130_fd_sc_hd__and2_1
X_4797_ _4797_/A vssd1 vssd1 vccd1 vccd1 _6463_/D sky130_fd_sc_hd__clkbuf_1
X_6536_ _6546_/CLK _6536_/D vssd1 vssd1 vccd1 vccd1 _6536_/Q sky130_fd_sc_hd__dfxtp_1
X_3748_ _3718_/X _3716_/C _3746_/X _5001_/A vssd1 vssd1 vccd1 vccd1 _3749_/B sky130_fd_sc_hd__a31o_1
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3679_ _3679_/A _3679_/B _3679_/C vssd1 vssd1 vccd1 vccd1 _3679_/X sky130_fd_sc_hd__and3_1
X_6467_ _6763_/CLK _6467_/D vssd1 vssd1 vccd1 vccd1 _6467_/Q sky130_fd_sc_hd__dfxtp_1
X_5418_ _3865_/A _3639_/A _5431_/S vssd1 vssd1 vccd1 vccd1 _5419_/B sky130_fd_sc_hd__mux2_1
X_6398_ _6789_/CLK _6398_/D vssd1 vssd1 vccd1 vccd1 _6398_/Q sky130_fd_sc_hd__dfxtp_1
X_5349_ _6626_/Q _5372_/B vssd1 vssd1 vccd1 vccd1 _5350_/A sky130_fd_sc_hd__and2_1
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6873__133 vssd1 vssd1 vccd1 vccd1 _6873__133/HI _6982_/A sky130_fd_sc_hd__conb_1
XFILLER_24_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _6373_/Q _4722_/B vssd1 vssd1 vccd1 vccd1 _4721_/A sky130_fd_sc_hd__and2_1
XFILLER_42_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4651_ _6334_/Q _4655_/B vssd1 vssd1 vccd1 vccd1 _4652_/A sky130_fd_sc_hd__and2_1
X_3602_ _3727_/A _3727_/B _3720_/C _3645_/B vssd1 vssd1 vccd1 vccd1 _3660_/A sky130_fd_sc_hd__nand4_2
Xinput31 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _3325_/D sky130_fd_sc_hd__buf_2
Xinput20 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _3333_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4582_ _4602_/B _4582_/B vssd1 vssd1 vccd1 vccd1 _4583_/B sky130_fd_sc_hd__xnor2_1
Xinput53 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 _4909_/B sky130_fd_sc_hd__clkbuf_4
Xinput42 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_4
Xinput64 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_4
X_6321_ _6528_/CLK _6321_/D vssd1 vssd1 vccd1 vccd1 _6321_/Q sky130_fd_sc_hd__dfxtp_1
X_3533_ _3569_/C _3533_/B vssd1 vssd1 vccd1 vccd1 _3538_/A sky130_fd_sc_hd__or2_1
XFILLER_115_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3464_ _3486_/A vssd1 vssd1 vccd1 vccd1 _3473_/S sky130_fd_sc_hd__clkbuf_2
X_6252_ _6805_/Q _6247_/X _6251_/Y _6235_/X vssd1 vssd1 vccd1 vccd1 _6805_/D sky130_fd_sc_hd__o211a_1
X_5203_ _5203_/A vssd1 vssd1 vccd1 vccd1 _6584_/D sky130_fd_sc_hd__clkbuf_1
X_6183_ _6783_/Q _6169_/A _6182_/X _6178_/X vssd1 vssd1 vccd1 vccd1 _6783_/D sky130_fd_sc_hd__o211a_1
X_3395_ _6293_/Q _3396_/C _3394_/Y _3398_/B vssd1 vssd1 vccd1 vccd1 _6293_/D sky130_fd_sc_hd__o211a_1
XFILLER_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5134_ _5119_/X _5133_/X _5115_/X vssd1 vssd1 vccd1 vccd1 _5135_/C sky130_fd_sc_hd__a21o_1
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _5077_/A _5065_/B vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__or2_1
X_4016_ _4033_/C _4016_/B vssd1 vssd1 vccd1 vccd1 _4017_/B sky130_fd_sc_hd__xnor2_2
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6857__117 vssd1 vssd1 vccd1 vccd1 _6857__117/HI _6966_/A sky130_fd_sc_hd__conb_1
XFILLER_92_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5967_ _6058_/A vssd1 vssd1 vccd1 vccd1 _6023_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4918_ _4918_/A vssd1 vssd1 vccd1 vccd1 _6527_/D sky130_fd_sc_hd__clkbuf_1
X_5898_ _6481_/Q _5964_/D _5914_/C vssd1 vssd1 vccd1 vccd1 _5898_/X sky130_fd_sc_hd__and3_1
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4849_ _4849_/A vssd1 vssd1 vccd1 vccd1 _6486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6519_ _6531_/CLK _6519_/D vssd1 vssd1 vccd1 vccd1 _6519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ input1/X vssd1 vssd1 vccd1 vccd1 _3305_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6836__96 vssd1 vssd1 vccd1 vccd1 _6836__96/HI _6945_/A sky130_fd_sc_hd__conb_1
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5821_ _5581_/X _5819_/X _5842_/S vssd1 vssd1 vccd1 vccd1 _5821_/X sky130_fd_sc_hd__mux2_1
X_5752_ _5630_/X _5751_/X _5757_/S vssd1 vssd1 vccd1 vccd1 _5752_/X sky130_fd_sc_hd__mux2_1
X_4703_ _6365_/Q _4711_/B vssd1 vssd1 vccd1 vccd1 _4704_/A sky130_fd_sc_hd__and2_1
X_5683_ _5882_/A _5882_/B vssd1 vssd1 vccd1 vccd1 _6059_/A sky130_fd_sc_hd__nand2_2
X_4634_ _4634_/A vssd1 vssd1 vccd1 vccd1 _4634_/Y sky130_fd_sc_hd__inv_2
X_4565_ _4613_/B _4565_/B vssd1 vssd1 vccd1 vccd1 _4615_/B sky130_fd_sc_hd__or2_1
X_6304_ _6504_/CLK _6304_/D vssd1 vssd1 vccd1 vccd1 _6304_/Q sky130_fd_sc_hd__dfxtp_1
X_3516_ _6649_/Q _6648_/Q _3534_/B _3516_/D vssd1 vssd1 vccd1 vccd1 _3539_/A sky130_fd_sc_hd__and4_1
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4496_ _4597_/B vssd1 vssd1 vccd1 vccd1 _4637_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6235_ _6255_/A vssd1 vssd1 vccd1 vccd1 _6235_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3447_ _3881_/A _6507_/Q _3451_/S vssd1 vssd1 vccd1 vccd1 _3448_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3378_ _4259_/A vssd1 vssd1 vccd1 vccd1 _5193_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6776_/Q _6156_/X _6164_/X _6165_/X vssd1 vssd1 vccd1 vccd1 _6776_/D sky130_fd_sc_hd__o211a_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5117_ _6908_/A _5041_/A _5116_/X _5100_/X vssd1 vssd1 vccd1 vccd1 _6570_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6468_/Q _6081_/X _6096_/X _6087_/X _6484_/Q vssd1 vssd1 vccd1 vccd1 _6097_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5048_ _5113_/A vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_85_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6999_ _6999_/A _3307_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
XFILLER_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4350_ _4350_/A _4350_/B vssd1 vssd1 vccd1 vccd1 _4350_/Y sky130_fd_sc_hd__nand2_1
X_3301_ _3304_/A vssd1 vssd1 vccd1 vccd1 _3301_/Y sky130_fd_sc_hd__inv_2
X_4281_ _4433_/C vssd1 vssd1 vccd1 vccd1 _4373_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3232_ _3250_/A vssd1 vssd1 vccd1 vccd1 _3237_/A sky130_fd_sc_hd__buf_12
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6020_ _6744_/Q _6011_/X _6019_/X _5999_/X vssd1 vssd1 vccd1 vccd1 _6744_/D sky130_fd_sc_hd__o211a_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6922_ _6922_/A _3215_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__ebufn_8
XFILLER_81_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5804_ _6481_/Q _5787_/X _5803_/X _5777_/X _5788_/X vssd1 vssd1 vccd1 vccd1 _5804_/X
+ sky130_fd_sc_hd__a221o_1
X_6784_ _6799_/CLK _6784_/D vssd1 vssd1 vccd1 vccd1 _6784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3996_ _3944_/A _4114_/C _4153_/C _3944_/B vssd1 vssd1 vccd1 vccd1 _4000_/C sky130_fd_sc_hd__a22o_1
X_5735_ _5735_/A vssd1 vssd1 vccd1 vccd1 _5735_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5666_ _6686_/Q _5650_/X _5663_/X _5665_/X _5640_/X vssd1 vssd1 vccd1 vccd1 _6686_/D
+ sky130_fd_sc_hd__o221a_1
X_4617_ _4614_/X _4615_/X _4612_/Y vssd1 vssd1 vccd1 vccd1 _4618_/B sky130_fd_sc_hd__a21o_1
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5597_ _5593_/X _5582_/X _5571_/X _5596_/X vssd1 vssd1 vccd1 vccd1 _5597_/X sky130_fd_sc_hd__o211a_1
X_4548_ _6671_/Q vssd1 vssd1 vccd1 vccd1 _4622_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4479_ _4543_/A _4479_/B _4576_/C _6379_/Q vssd1 vssd1 vccd1 vccd1 _4480_/B sky130_fd_sc_hd__and4_1
X_6218_ _6280_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6218_/X sky130_fd_sc_hd__or2_1
XFILLER_58_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6149_ _6237_/A _6154_/B vssd1 vssd1 vccd1 vccd1 _6149_/X sky130_fd_sc_hd__or2_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3850_ _3850_/A _3881_/A _3850_/C vssd1 vssd1 vccd1 vccd1 _3853_/A sky130_fd_sc_hd__and3_1
X_3781_ _5441_/A vssd1 vssd1 vccd1 vccd1 _3781_/X sky130_fd_sc_hd__buf_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5520_ _6478_/Q _5638_/A _6056_/C _5519_/X vssd1 vssd1 vccd1 vccd1 _5520_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5451_ _5469_/A vssd1 vssd1 vccd1 vccd1 _5466_/S sky130_fd_sc_hd__buf_2
X_5382_ _6643_/Q _6642_/Q _6641_/Q vssd1 vssd1 vccd1 vccd1 _5668_/B sky130_fd_sc_hd__nor3_4
X_4402_ _4429_/A _4450_/B _4429_/C vssd1 vssd1 vccd1 vccd1 _4404_/B sky130_fd_sc_hd__nand3_1
XFILLER_99_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4333_ _4333_/A _4333_/B vssd1 vssd1 vccd1 vccd1 _4340_/A sky130_fd_sc_hd__nand2_1
XFILLER_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4264_ _4264_/A _4270_/B vssd1 vssd1 vccd1 vccd1 _4265_/A sky130_fd_sc_hd__and2_1
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3215_ _3218_/A vssd1 vssd1 vccd1 vccd1 _3215_/Y sky130_fd_sc_hd__inv_2
X_6003_ _6003_/A vssd1 vssd1 vccd1 vccd1 _6003_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4195_ _4218_/B _4195_/B _4220_/D vssd1 vssd1 vccd1 vccd1 _4195_/X sky130_fd_sc_hd__or3_1
XFILLER_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6905_ _6905_/A _3193_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__ebufn_8
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6820__80 vssd1 vssd1 vccd1 vccd1 _6820__80/HI _6929_/A sky130_fd_sc_hd__conb_1
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6767_ _6799_/CLK _6767_/D vssd1 vssd1 vccd1 vccd1 _6767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3979_ _3973_/X _3977_/X _4151_/A _3979_/D vssd1 vssd1 vccd1 vccd1 _4009_/A sky130_fd_sc_hd__and4bb_1
X_5718_ _5797_/A vssd1 vssd1 vccd1 vccd1 _5718_/X sky130_fd_sc_hd__clkbuf_2
X_6698_ _6809_/CLK _6698_/D vssd1 vssd1 vccd1 vccd1 _6698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5649_ _6684_/Q _5601_/X _5646_/X _5648_/X _5640_/X vssd1 vssd1 vccd1 vccd1 _6684_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4951_ _4950_/B _5118_/B _4950_/A vssd1 vssd1 vccd1 vccd1 _4952_/C sky130_fd_sc_hd__a21o_1
XFILLER_24_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4882_ _6505_/Q _4880_/X _4881_/X input63/X vssd1 vssd1 vccd1 vccd1 _6505_/D sky130_fd_sc_hd__a22o_1
X_3902_ _6352_/Q vssd1 vssd1 vccd1 vccd1 _3998_/C sky130_fd_sc_hd__clkbuf_2
X_6621_ _6799_/CLK _6621_/D vssd1 vssd1 vccd1 vccd1 _6621_/Q sky130_fd_sc_hd__dfxtp_1
X_3833_ _3822_/B _3833_/B vssd1 vssd1 vccd1 vccd1 _3843_/A sky130_fd_sc_hd__and2b_1
X_6552_ _6554_/CLK _6552_/D vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfxtp_2
X_3764_ _3764_/A _3764_/B vssd1 vssd1 vccd1 vccd1 _3766_/A sky130_fd_sc_hd__xnor2_1
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5503_ _5535_/A vssd1 vssd1 vccd1 vccd1 _6040_/A sky130_fd_sc_hd__clkbuf_2
X_6483_ _6763_/CLK _6483_/D vssd1 vssd1 vccd1 vccd1 _6483_/Q sky130_fd_sc_hd__dfxtp_4
X_3695_ _3656_/A _3656_/C _3656_/B vssd1 vssd1 vccd1 vccd1 _3696_/C sky130_fd_sc_hd__a21bo_1
X_5434_ _5469_/A vssd1 vssd1 vccd1 vccd1 _5448_/S sky130_fd_sc_hd__buf_2
XFILLER_99_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5365_ _5363_/Y _5364_/X _4352_/X vssd1 vssd1 vccd1 vccd1 _6629_/D sky130_fd_sc_hd__o21ai_1
X_5296_ _5374_/A vssd1 vssd1 vccd1 vccd1 _5305_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4316_ _6665_/Q _4333_/B _4354_/B _6664_/Q vssd1 vssd1 vccd1 vccd1 _4316_/X sky130_fd_sc_hd__a22o_1
X_4247_ _4247_/A _4247_/B _4247_/C vssd1 vssd1 vccd1 vccd1 _4249_/A sky130_fd_sc_hd__and3_1
X_4178_ _6663_/Q vssd1 vssd1 vccd1 vccd1 _4227_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3480_ _6318_/Q _6522_/Q _3484_/S vssd1 vssd1 vccd1 vccd1 _3481_/A sky130_fd_sc_hd__mux2_1
X_5150_ _5181_/A vssd1 vssd1 vccd1 vccd1 _5150_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5081_ _5081_/A vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4101_ _4101_/A vssd1 vssd1 vccd1 vccd1 _4230_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4032_ _4230_/C vssd1 vssd1 vccd1 vccd1 _4273_/A sky130_fd_sc_hd__buf_2
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5983_ _6737_/Q _5946_/X _5982_/X _5959_/X vssd1 vssd1 vccd1 vccd1 _6737_/D sky130_fd_sc_hd__o211a_1
XFILLER_52_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4934_ _5188_/A vssd1 vssd1 vccd1 vccd1 _4950_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_52_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_12 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _3313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4865_ _4865_/A vssd1 vssd1 vccd1 vccd1 _6493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6604_ _6667_/CLK _6604_/D vssd1 vssd1 vccd1 vccd1 _6604_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_34 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3816_ _3787_/A _5214_/A _3796_/B _3815_/X vssd1 vssd1 vccd1 vccd1 _3818_/B sky130_fd_sc_hd__a31oi_1
XFILLER_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4796_ _6415_/Q _4800_/B vssd1 vssd1 vccd1 vccd1 _4797_/A sky130_fd_sc_hd__and2_1
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6535_ _6570_/CLK _6535_/D vssd1 vssd1 vccd1 vccd1 _6535_/Q sky130_fd_sc_hd__dfxtp_1
X_3747_ _3718_/X _3716_/C _3746_/X vssd1 vssd1 vccd1 vccd1 _3749_/A sky130_fd_sc_hd__a21oi_1
X_3678_ _3638_/X _3639_/X _3667_/A _3668_/Y vssd1 vssd1 vccd1 vccd1 _3678_/Y sky130_fd_sc_hd__o211ai_2
X_6466_ _6763_/CLK _6466_/D vssd1 vssd1 vccd1 vccd1 _6466_/Q sky130_fd_sc_hd__dfxtp_1
X_6397_ _6795_/CLK _6397_/D vssd1 vssd1 vccd1 vccd1 _6397_/Q sky130_fd_sc_hd__dfxtp_1
X_5417_ _5496_/S vssd1 vssd1 vccd1 vccd1 _5431_/S sky130_fd_sc_hd__buf_2
X_5348_ _5374_/A vssd1 vssd1 vccd1 vccd1 _5372_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5279_ _5279_/A vssd1 vssd1 vccd1 vccd1 _6604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4650_ _4647_/A _4649_/X _4255_/X vssd1 vssd1 vccd1 vccd1 _6397_/D sky130_fd_sc_hd__o21a_1
Xinput21 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _3333_/D sky130_fd_sc_hd__clkbuf_2
X_3601_ _6299_/Q vssd1 vssd1 vccd1 vccd1 _3720_/C sky130_fd_sc_hd__clkbuf_2
Xinput10 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 _3331_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_30_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput32 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _3325_/C sky130_fd_sc_hd__clkbuf_2
Xinput54 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 _4912_/B sky130_fd_sc_hd__clkbuf_4
X_6320_ _6531_/CLK _6320_/D vssd1 vssd1 vccd1 vccd1 _6320_/Q sky130_fd_sc_hd__dfxtp_1
X_4581_ _4552_/A _4551_/A _4551_/B vssd1 vssd1 vccd1 vccd1 _4582_/B sky130_fd_sc_hd__o21ba_1
Xinput43 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_4
Xinput65 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_6
XFILLER_115_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3532_ _3729_/A _3516_/D _3578_/B _3755_/B vssd1 vssd1 vccd1 vccd1 _3533_/B sky130_fd_sc_hd__a22oi_1
X_3463_ _3463_/A vssd1 vssd1 vccd1 vccd1 _6310_/D sky130_fd_sc_hd__clkbuf_1
X_6251_ _6248_/X _6250_/Y _6244_/X vssd1 vssd1 vccd1 vccd1 _6251_/Y sky130_fd_sc_hd__o21ai_1
X_5202_ _5243_/A _5202_/B _5202_/C vssd1 vssd1 vccd1 vccd1 _5203_/A sky130_fd_sc_hd__and3_1
X_6182_ _6286_/A _6182_/B vssd1 vssd1 vccd1 vccd1 _6182_/X sky130_fd_sc_hd__or2_1
X_3394_ _6293_/Q _3396_/C vssd1 vssd1 vccd1 vccd1 _3394_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5133_ _6690_/Q _6722_/Q _6754_/Q _6786_/Q _5126_/X _4950_/A vssd1 vssd1 vccd1 vccd1
+ _5133_/X sky130_fd_sc_hd__mux4_2
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5064_ _6679_/Q _6711_/Q _6743_/Q _6775_/Q _5049_/X _5063_/X vssd1 vssd1 vccd1 vccd1
+ _5065_/B sky130_fd_sc_hd__mux4_1
X_4015_ _6657_/Q _4151_/B vssd1 vssd1 vccd1 vccd1 _4016_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5966_ _6622_/Q _6224_/C vssd1 vssd1 vccd1 vccd1 _6058_/A sky130_fd_sc_hd__and2_1
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4917_ _4916_/X _6527_/Q _4926_/S vssd1 vssd1 vccd1 vccd1 _4918_/A sky130_fd_sc_hd__mux2_1
X_5897_ _5552_/X _5889_/X _5891_/X _5874_/X _6723_/Q vssd1 vssd1 vccd1 vccd1 _5897_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_33_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4848_ _6438_/Q _4856_/B vssd1 vssd1 vccd1 vccd1 _4849_/A sky130_fd_sc_hd__and2_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _4779_/A vssd1 vssd1 vccd1 vccd1 _6455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6518_ _6531_/CLK _6518_/D vssd1 vssd1 vccd1 vccd1 _6518_/Q sky130_fd_sc_hd__dfxtp_1
X_6449_ _6789_/CLK _6449_/D vssd1 vssd1 vccd1 vccd1 _6449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6840__100 vssd1 vssd1 vccd1 vccd1 _6840__100/HI _6949_/A sky130_fd_sc_hd__conb_1
XFILLER_48_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5820_ _5866_/S vssd1 vssd1 vccd1 vccd1 _5842_/S sky130_fd_sc_hd__clkbuf_2
X_5751_ _6699_/Q _5633_/X _5751_/S vssd1 vssd1 vccd1 vccd1 _5751_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4702_ _4735_/A vssd1 vssd1 vccd1 vccd1 _4711_/B sky130_fd_sc_hd__clkbuf_1
X_5682_ _6688_/Q _5508_/X _5764_/S vssd1 vssd1 vccd1 vccd1 _5682_/X sky130_fd_sc_hd__mux2_1
X_4633_ _4614_/X _4615_/X _4630_/Y _4612_/Y vssd1 vssd1 vccd1 vccd1 _4633_/X sky130_fd_sc_hd__a211o_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4564_ _4613_/A _4563_/B _4563_/C vssd1 vssd1 vccd1 vccd1 _4565_/B sky130_fd_sc_hd__o21a_1
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6303_ _6509_/CLK _6303_/D vssd1 vssd1 vccd1 vccd1 _6303_/Q sky130_fd_sc_hd__dfxtp_1
X_3515_ _3515_/A vssd1 vssd1 vccd1 vccd1 _6335_/D sky130_fd_sc_hd__clkbuf_1
X_4495_ _4492_/X _4493_/Y _4468_/X _4455_/X vssd1 vssd1 vccd1 vccd1 _4502_/C sky130_fd_sc_hd__a211o_1
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6234_ _6227_/X _6233_/Y _6230_/X vssd1 vssd1 vccd1 vccd1 _6234_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3446_ _5214_/A vssd1 vssd1 vccd1 vccd1 _3881_/A sky130_fd_sc_hd__clkbuf_2
X_3377_ _3377_/A vssd1 vssd1 vccd1 vccd1 _4259_/A sky130_fd_sc_hd__buf_4
XFILLER_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6165_ _6178_/A vssd1 vssd1 vccd1 vccd1 _6165_/X sky130_fd_sc_hd__buf_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5116_ _5081_/A _5113_/X _5114_/X _5115_/X vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__a31o_1
XFILLER_85_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6096_ _6096_/A vssd1 vssd1 vccd1 vccd1 _6096_/X sky130_fd_sc_hd__clkbuf_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5047_ _5081_/A vssd1 vssd1 vccd1 vccd1 _5047_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6998_ _6998_/A _3306_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
XFILLER_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5949_ _6490_/Q _5957_/B _5957_/C vssd1 vssd1 vccd1 vccd1 _5949_/X sky130_fd_sc_hd__and3_1
XFILLER_40_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3300_ _3304_/A vssd1 vssd1 vccd1 vccd1 _3300_/Y sky130_fd_sc_hd__inv_2
X_4280_ _6374_/Q vssd1 vssd1 vccd1 vccd1 _4433_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3231_ _3231_/A vssd1 vssd1 vccd1 vccd1 _3231_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6921_ _6921_/A _3214_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__ebufn_8
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5803_ _5552_/X _5802_/X _5814_/S vssd1 vssd1 vccd1 vccd1 _5803_/X sky130_fd_sc_hd__mux2_1
X_6783_ _6799_/CLK _6783_/D vssd1 vssd1 vccd1 vccd1 _6783_/Q sky130_fd_sc_hd__dfxtp_1
X_3995_ _3995_/A _3995_/B vssd1 vssd1 vccd1 vccd1 _4067_/A sky130_fd_sc_hd__nand2_1
X_5734_ _5734_/A vssd1 vssd1 vccd1 vccd1 _5734_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5665_ _6283_/A _5638_/X _5627_/X _5519_/X vssd1 vssd1 vccd1 vccd1 _5665_/X sky130_fd_sc_hd__a31o_1
X_4616_ _4612_/Y _4614_/X _4615_/X _3636_/A vssd1 vssd1 vccd1 vccd1 _4616_/X sky130_fd_sc_hd__a31o_1
X_5596_ _5624_/A _5596_/B vssd1 vssd1 vccd1 vccd1 _5596_/X sky130_fd_sc_hd__or2_1
X_4547_ _4547_/A _4547_/B vssd1 vssd1 vccd1 vccd1 _4552_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4478_ _4543_/A _4512_/B _4547_/B _4545_/B vssd1 vssd1 vccd1 vccd1 _4480_/A sky130_fd_sc_hd__a22oi_1
X_6217_ _6796_/Q _6207_/X _6215_/X _6216_/X vssd1 vssd1 vccd1 vccd1 _6796_/D sky130_fd_sc_hd__o211a_1
X_3429_ _6301_/Q vssd1 vssd1 vccd1 vccd1 _3789_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6148_ _6769_/Q _6142_/X _6147_/X _6051_/X vssd1 vssd1 vccd1 vccd1 _6769_/D sky130_fd_sc_hd__o211a_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6079_ _6079_/A vssd1 vssd1 vccd1 vccd1 _6754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3780_ _3828_/A _3828_/C _3779_/X vssd1 vssd1 vccd1 vccd1 _3780_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5450_ _5450_/A vssd1 vssd1 vccd1 vccd1 _6657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4401_ _4401_/A _4437_/A vssd1 vssd1 vccd1 vccd1 _4429_/C sky130_fd_sc_hd__nor2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5381_ _6647_/Q _6646_/Q _6645_/Q _6644_/Q vssd1 vssd1 vccd1 vccd1 _5383_/A sky130_fd_sc_hd__or4_1
XFILLER_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_4332_ _4332_/A _4332_/B vssd1 vssd1 vccd1 vccd1 _4342_/A sky130_fd_sc_hd__xnor2_1
XFILLER_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4263_ _4263_/A vssd1 vssd1 vccd1 vccd1 _6375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6002_ _6741_/Q _5570_/X _6017_/S vssd1 vssd1 vccd1 vccd1 _6002_/X sky130_fd_sc_hd__mux2_1
X_3214_ _3218_/A vssd1 vssd1 vccd1 vccd1 _3214_/Y sky130_fd_sc_hd__inv_2
X_4194_ _4218_/A _4194_/B vssd1 vssd1 vccd1 vccd1 _4220_/D sky130_fd_sc_hd__xor2_1
XFILLER_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6904_ _6904_/A _3192_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__ebufn_8
XFILLER_54_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6766_ _6795_/CLK _6766_/D vssd1 vssd1 vccd1 vccd1 _6766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3978_ _6661_/Q vssd1 vssd1 vccd1 vccd1 _4151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5717_ _6692_/Q _5650_/X _5715_/X _5716_/X _5707_/X vssd1 vssd1 vccd1 vccd1 _6692_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6697_ _6809_/CLK _6697_/D vssd1 vssd1 vccd1 vccd1 _6697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5648_ _6277_/A _5638_/X _5627_/X _5616_/X vssd1 vssd1 vccd1 vccd1 _5648_/X sky130_fd_sc_hd__a31o_1
XFILLER_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5579_ _6250_/A _5534_/X _5578_/X _5567_/X vssd1 vssd1 vccd1 vccd1 _5579_/X sky130_fd_sc_hd__a31o_1
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput8 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4950_ _4950_/A _4950_/B _5118_/B vssd1 vssd1 vccd1 vccd1 _4950_/X sky130_fd_sc_hd__and3_1
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3901_ _5162_/A vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__buf_2
X_4881_ _4895_/A vssd1 vssd1 vccd1 vccd1 _4881_/X sky130_fd_sc_hd__clkbuf_2
X_6620_ _6799_/CLK _6620_/D vssd1 vssd1 vccd1 vccd1 _6620_/Q sky130_fd_sc_hd__dfxtp_1
X_3832_ _3832_/A vssd1 vssd1 vccd1 vccd1 _6346_/D sky130_fd_sc_hd__clkbuf_1
X_6551_ _6551_/CLK _6551_/D vssd1 vssd1 vccd1 vccd1 _6551_/Q sky130_fd_sc_hd__dfxtp_1
X_5502_ _5880_/A _5502_/B _5775_/B vssd1 vssd1 vccd1 vccd1 _5535_/A sky130_fd_sc_hd__nor3_1
X_3763_ _3763_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3764_/B sky130_fd_sc_hd__nor2_1
X_6482_ _6763_/CLK _6482_/D vssd1 vssd1 vccd1 vccd1 _6482_/Q sky130_fd_sc_hd__dfxtp_4
X_3694_ _3694_/A _3694_/B _3694_/C vssd1 vssd1 vccd1 vccd1 _3696_/B sky130_fd_sc_hd__nand3_1
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5433_ _5433_/A vssd1 vssd1 vccd1 vccd1 _6652_/D sky130_fd_sc_hd__clkbuf_1
X_5364_ _6629_/Q _5364_/B vssd1 vssd1 vccd1 vccd1 _5364_/X sky130_fd_sc_hd__and2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4315_ _6665_/Q _6664_/Q _4333_/B vssd1 vssd1 vccd1 vccd1 _4315_/X sky130_fd_sc_hd__and3_1
X_5295_ _5295_/A vssd1 vssd1 vccd1 vccd1 _6611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4246_ _4246_/A vssd1 vssd1 vccd1 vccd1 _4247_/C sky130_fd_sc_hd__inv_2
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4177_ _4177_/A _4230_/D vssd1 vssd1 vccd1 vccd1 _4187_/A sky130_fd_sc_hd__nand2_2
XFILLER_67_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6749_ _6532_/Q _6749_/D vssd1 vssd1 vccd1 vccd1 _6749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5080_ _6902_/A _5075_/X _5079_/X _5068_/X vssd1 vssd1 vccd1 vccd1 _6564_/D sky130_fd_sc_hd__o211a_1
X_4100_ _4097_/X _4098_/Y _4074_/X _4062_/X vssd1 vssd1 vccd1 vccd1 _4106_/C sky130_fd_sc_hd__a211o_1
XFILLER_84_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4031_ _4058_/B vssd1 vssd1 vccd1 vccd1 _4230_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_65_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5982_ _5969_/X _5980_/X _5981_/X vssd1 vssd1 vccd1 vccd1 _5982_/X sky130_fd_sc_hd__a21o_1
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4933_ _6533_/Q vssd1 vssd1 vccd1 vccd1 _5188_/A sky130_fd_sc_hd__buf_2
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4864_ _6445_/Q _4959_/B vssd1 vssd1 vccd1 vccd1 _4865_/A sky130_fd_sc_hd__and2_1
XANTENNA_13 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6603_ _6667_/CLK _6603_/D vssd1 vssd1 vccd1 vccd1 _6603_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_24 _3231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3815_ _3795_/B _3815_/B vssd1 vssd1 vccd1 vccd1 _3815_/X sky130_fd_sc_hd__and2b_1
XANTENNA_35 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4795_ _4795_/A vssd1 vssd1 vccd1 vccd1 _6462_/D sky130_fd_sc_hd__clkbuf_1
X_6534_ _6570_/CLK _6534_/D vssd1 vssd1 vccd1 vccd1 _6534_/Q sky130_fd_sc_hd__dfxtp_1
X_3746_ _3778_/C _3745_/Y vssd1 vssd1 vccd1 vccd1 _3746_/X sky130_fd_sc_hd__or2b_1
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6465_ _6809_/CLK _6465_/D vssd1 vssd1 vccd1 vccd1 _6465_/Q sky130_fd_sc_hd__dfxtp_1
X_5416_ _5469_/A vssd1 vssd1 vccd1 vccd1 _5496_/S sky130_fd_sc_hd__buf_2
X_3677_ _4990_/A _3677_/B vssd1 vssd1 vccd1 vccd1 _6341_/D sky130_fd_sc_hd__nor2_1
X_6396_ _6795_/CLK _6396_/D vssd1 vssd1 vccd1 vccd1 _6396_/Q sky130_fd_sc_hd__dfxtp_1
X_5347_ _5347_/A vssd1 vssd1 vccd1 vccd1 _6625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5278_ _6604_/Q _5282_/B vssd1 vssd1 vccd1 vccd1 _5279_/A sky130_fd_sc_hd__and2_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4229_ _4242_/A _4230_/C _4230_/D _4241_/A vssd1 vssd1 vccd1 vccd1 _4231_/A sky130_fd_sc_hd__a22o_1
XFILLER_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4580_ _4580_/A _4600_/B vssd1 vssd1 vccd1 vccd1 _4602_/B sky130_fd_sc_hd__nor2_1
Xinput22 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _3333_/C sky130_fd_sc_hd__clkbuf_2
X_3600_ _6651_/Q _6299_/Q _3645_/B _6652_/Q vssd1 vssd1 vccd1 vccd1 _3605_/C sky130_fd_sc_hd__a22o_1
Xinput11 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _3331_/A sky130_fd_sc_hd__buf_2
XFILLER_30_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput55 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 _4916_/B sky130_fd_sc_hd__clkbuf_2
Xinput44 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_4
Xinput33 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _3327_/B sky130_fd_sc_hd__buf_4
X_3531_ _3755_/B _3650_/A _3556_/C _3578_/B vssd1 vssd1 vccd1 vccd1 _3569_/C sky130_fd_sc_hd__and4_1
Xinput66 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3462_ _6310_/Q _6514_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _3463_/A sky130_fd_sc_hd__mux2_1
X_6250_ _6250_/A _6263_/B vssd1 vssd1 vccd1 vccd1 _6250_/Y sky130_fd_sc_hd__nand2_1
X_3393_ _3393_/A vssd1 vssd1 vccd1 vccd1 _6292_/D sky130_fd_sc_hd__clkbuf_1
X_5201_ _5181_/X _5200_/X _5176_/X vssd1 vssd1 vccd1 vccd1 _5202_/C sky130_fd_sc_hd__a21o_1
X_6181_ _6782_/Q _6169_/X _6180_/X _6178_/X vssd1 vssd1 vccd1 vccd1 _6782_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5132_ _6911_/A _5149_/B vssd1 vssd1 vccd1 vccd1 _5135_/B sky130_fd_sc_hd__or2_1
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5063_ _5169_/A vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__clkbuf_2
X_4014_ _4123_/A _3998_/D _3977_/D _3972_/X vssd1 vssd1 vccd1 vccd1 _4033_/C sky130_fd_sc_hd__a31o_1
XFILLER_92_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5965_ _5963_/X _5964_/X _5331_/X vssd1 vssd1 vccd1 vccd1 _6735_/D sky130_fd_sc_hd__o21a_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4916_ _4919_/A _4916_/B vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__and2_1
X_5896_ _6722_/Q _5888_/X _5895_/X _5863_/X vssd1 vssd1 vccd1 vccd1 _6722_/D sky130_fd_sc_hd__o211a_1
X_4847_ _4847_/A vssd1 vssd1 vccd1 vccd1 _4856_/B sky130_fd_sc_hd__clkbuf_1
X_4778_ _6407_/Q _4778_/B vssd1 vssd1 vccd1 vccd1 _4779_/A sky130_fd_sc_hd__and2_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6517_ _6528_/CLK _6517_/D vssd1 vssd1 vccd1 vccd1 _6517_/Q sky130_fd_sc_hd__dfxtp_1
X_3729_ _3729_/A _6303_/Q vssd1 vssd1 vccd1 vccd1 _3751_/B sky130_fd_sc_hd__nand2_1
X_6448_ _6789_/CLK _6448_/D vssd1 vssd1 vccd1 vccd1 _6448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6379_ _6795_/CLK _6379_/D vssd1 vssd1 vccd1 vccd1 _6379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5750_ _6698_/Q _5380_/X _5748_/X _5749_/X _5707_/X vssd1 vssd1 vccd1 vccd1 _6698_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _5770_/S vssd1 vssd1 vccd1 vccd1 _5764_/S sky130_fd_sc_hd__buf_2
X_4701_ _4701_/A vssd1 vssd1 vccd1 vccd1 _6420_/D sky130_fd_sc_hd__clkbuf_1
X_4632_ _4634_/A _4618_/B _4630_/Y _4631_/Y _3633_/X vssd1 vssd1 vccd1 vccd1 _6395_/D
+ sky130_fd_sc_hd__a311oi_1
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4563_ _4613_/A _4563_/B _4563_/C vssd1 vssd1 vccd1 vccd1 _4613_/B sky130_fd_sc_hd__nor3_1
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4494_ _4468_/X _4455_/X _4492_/X _4493_/Y vssd1 vssd1 vccd1 vccd1 _4502_/B sky130_fd_sc_hd__o211ai_2
X_6302_ _6509_/CLK _6302_/D vssd1 vssd1 vccd1 vccd1 _6302_/Q sky130_fd_sc_hd__dfxtp_1
X_3514_ _3899_/A _3514_/B _3526_/A vssd1 vssd1 vccd1 vccd1 _3515_/A sky130_fd_sc_hd__and3_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3445_ _3810_/B vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__clkbuf_2
X_6233_ _6233_/A _6243_/B vssd1 vssd1 vccd1 vccd1 _6233_/Y sky130_fd_sc_hd__nand2_1
X_6863__123 vssd1 vssd1 vccd1 vccd1 _6863__123/HI _6972_/A sky130_fd_sc_hd__conb_1
X_3376_ _6289_/Q _6330_/D vssd1 vssd1 vccd1 vccd1 _6289_/D sky130_fd_sc_hd__nor2_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6260_/A _6167_/B vssd1 vssd1 vccd1 vccd1 _6164_/X sky130_fd_sc_hd__or2_1
X_5115_ _5176_/A vssd1 vssd1 vccd1 vccd1 _5115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6827__87 vssd1 vssd1 vccd1 vccd1 _6827__87/HI _6936_/A sky130_fd_sc_hd__conb_1
X_6095_ _6095_/A vssd1 vssd1 vccd1 vccd1 _6757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5046_ _6897_/A _5041_/X _5045_/X _5034_/X vssd1 vssd1 vccd1 vccd1 _6559_/D sky130_fd_sc_hd__o211a_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6997_ _6997_/A _3304_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
X_5948_ _5642_/X _5947_/X _5920_/A _5961_/B _6732_/Q vssd1 vssd1 vccd1 vccd1 _5948_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5879_ _5879_/A _5879_/B vssd1 vssd1 vccd1 vccd1 _6720_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6528_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6847__107 vssd1 vssd1 vccd1 vccd1 _6847__107/HI _6956_/A sky130_fd_sc_hd__conb_1
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3231_/A vssd1 vssd1 vccd1 vccd1 _3230_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6920_ _6920_/A _3212_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__ebufn_8
XFILLER_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5802_ _6707_/Q _5553_/X _5813_/S vssd1 vssd1 vccd1 vccd1 _5802_/X sky130_fd_sc_hd__mux2_1
X_6782_ _6532_/Q _6782_/D vssd1 vssd1 vccd1 vccd1 _6782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3994_ _3994_/A vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__inv_2
X_5733_ _6695_/Q _5718_/X _5732_/X _5690_/X vssd1 vssd1 vccd1 vccd1 _6695_/D sky130_fd_sc_hd__o211a_1
X_5664_ _6492_/Q vssd1 vssd1 vccd1 vccd1 _6283_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4615_ _4615_/A _4615_/B _4615_/C _4615_/D vssd1 vssd1 vccd1 vccd1 _4615_/X sky130_fd_sc_hd__or4_1
X_5595_ _6679_/Q _5594_/X _5612_/S vssd1 vssd1 vccd1 vccd1 _5596_/B sky130_fd_sc_hd__mux2_1
X_4546_ _4546_/A _4588_/A vssd1 vssd1 vccd1 vccd1 _4584_/A sky130_fd_sc_hd__or2_1
XFILLER_104_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4477_ _4477_/A _6380_/Q vssd1 vssd1 vccd1 vccd1 _4481_/A sky130_fd_sc_hd__nand2_1
X_3428_ _3428_/A vssd1 vssd1 vccd1 vccd1 _6300_/D sky130_fd_sc_hd__clkbuf_1
X_6216_ _6255_/A vssd1 vssd1 vccd1 vccd1 _6216_/X sky130_fd_sc_hd__buf_4
XFILLER_100_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3359_ _3357_/X _3358_/X _3340_/X vssd1 vssd1 vccd1 vccd1 _6329_/D sky130_fd_sc_hd__o21a_1
X_6147_ _6233_/A _6154_/B vssd1 vssd1 vccd1 vccd1 _6147_/X sky130_fd_sc_hd__or2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6078_ _6084_/A _6078_/B vssd1 vssd1 vccd1 vccd1 _6079_/A sky130_fd_sc_hd__and2_1
XFILLER_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5029_ _5169_/A vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4400_ _4576_/B _6669_/Q _4433_/C _4400_/D vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__and4_1
X_5380_ _5650_/A vssd1 vssd1 vccd1 vccd1 _5380_/X sky130_fd_sc_hd__buf_2
X_4331_ _4407_/A _4388_/B vssd1 vssd1 vccd1 vccd1 _4332_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4262_ _4262_/A _4270_/B vssd1 vssd1 vccd1 vccd1 _4263_/A sky130_fd_sc_hd__and2_1
X_3213_ _3219_/A vssd1 vssd1 vccd1 vccd1 _3218_/A sky130_fd_sc_hd__buf_6
XFILLER_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6001_ _6029_/A vssd1 vssd1 vccd1 vccd1 _6001_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4193_ _4198_/A _4198_/B vssd1 vssd1 vccd1 vccd1 _4194_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6903_ _6903_/A _3191_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__ebufn_8
XFILLER_35_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6765_ _6795_/CLK _6765_/D vssd1 vssd1 vccd1 vccd1 _6765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3977_ _3972_/X _3998_/D _6658_/Q _3977_/D vssd1 vssd1 vccd1 vccd1 _3977_/X sky130_fd_sc_hd__and4b_1
XFILLER_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5716_ _6243_/A _5704_/X _5705_/X vssd1 vssd1 vccd1 vccd1 _5716_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6696_ _6809_/CLK _6696_/D vssd1 vssd1 vccd1 vccd1 _6696_/Q sky130_fd_sc_hd__dfxtp_1
X_5647_ _6490_/Q vssd1 vssd1 vccd1 vccd1 _6277_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_123_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5578_ _6269_/A vssd1 vssd1 vccd1 vccd1 _5578_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4529_ _4493_/B _4493_/Y _4527_/Y _4528_/X vssd1 vssd1 vccd1 vccd1 _4531_/B sky130_fd_sc_hd__a211o_1
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4880_ _4910_/S vssd1 vssd1 vccd1 vccd1 _4880_/X sky130_fd_sc_hd__clkbuf_2
X_3900_ _3900_/A vssd1 vssd1 vccd1 vccd1 _6359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3831_ _3829_/X _3831_/B vssd1 vssd1 vccd1 vccd1 _3832_/A sky130_fd_sc_hd__and2b_1
X_6550_ _6551_/CLK _6550_/D vssd1 vssd1 vccd1 vccd1 _6550_/Q sky130_fd_sc_hd__dfxtp_1
X_3762_ _3789_/A _3789_/B _3789_/D _3762_/D vssd1 vssd1 vccd1 vccd1 _3763_/B sky130_fd_sc_hd__and4_1
X_5501_ _5922_/A vssd1 vssd1 vccd1 vccd1 _5957_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6481_ _6763_/CLK _6481_/D vssd1 vssd1 vccd1 vccd1 _6481_/Q sky130_fd_sc_hd__dfxtp_4
X_3693_ _3694_/B _3694_/C _3694_/A vssd1 vssd1 vccd1 vccd1 _3696_/A sky130_fd_sc_hd__a21o_1
X_5432_ _5439_/A _5432_/B vssd1 vssd1 vccd1 vccd1 _5433_/A sky130_fd_sc_hd__and2_1
X_5363_ _6629_/Q _5364_/B vssd1 vssd1 vccd1 vccd1 _5363_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4314_ _4371_/B vssd1 vssd1 vccd1 vccd1 _4354_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5294_ _6611_/Q _5294_/B vssd1 vssd1 vccd1 vccd1 _5295_/A sky130_fd_sc_hd__and2_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4245_ _4245_/A _4245_/B vssd1 vssd1 vccd1 vccd1 _4246_/A sky130_fd_sc_hd__xnor2_1
XFILLER_67_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4176_ _4176_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _4198_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6748_ _6532_/Q _6748_/D vssd1 vssd1 vccd1 vccd1 _6748_/Q sky130_fd_sc_hd__dfxtp_1
X_6679_ _6532_/Q _6679_/D vssd1 vssd1 vccd1 vccd1 _6679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4030_ _3986_/X _4028_/X _4029_/Y vssd1 vssd1 vccd1 vccd1 _6364_/D sky130_fd_sc_hd__o21a_1
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5981_ _6479_/Q _6056_/B _6056_/C _5976_/X vssd1 vssd1 vccd1 vccd1 _5981_/X sky130_fd_sc_hd__a31o_1
X_4932_ _6532_/Q _4931_/X _3398_/B vssd1 vssd1 vccd1 vccd1 _6532_/D sky130_fd_sc_hd__o21ba_1
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_14 _4912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6602_ _6667_/CLK _6602_/D vssd1 vssd1 vccd1 vccd1 _6602_/Q sky130_fd_sc_hd__dfxtp_1
X_4863_ _4863_/A vssd1 vssd1 vccd1 vccd1 _6492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_25 _4255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ _3851_/A _3814_/B vssd1 vssd1 vccd1 vccd1 _3818_/A sky130_fd_sc_hd__or2_1
XANTENNA_36 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4794_ _6414_/Q _4800_/B vssd1 vssd1 vccd1 vccd1 _4795_/A sky130_fd_sc_hd__and2_1
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6533_ _6558_/CLK _6533_/D vssd1 vssd1 vccd1 vccd1 _6533_/Q sky130_fd_sc_hd__dfxtp_4
X_3745_ _3745_/A _3745_/B _3745_/C vssd1 vssd1 vccd1 vccd1 _3745_/Y sky130_fd_sc_hd__nand3_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6464_ _6809_/CLK _6464_/D vssd1 vssd1 vccd1 vccd1 _6464_/Q sky130_fd_sc_hd__dfxtp_1
X_5415_ _5415_/A _6588_/Q _5238_/B vssd1 vssd1 vccd1 vccd1 _5469_/A sky130_fd_sc_hd__or3b_4
X_3676_ _3676_/A _3676_/B vssd1 vssd1 vccd1 vccd1 _3677_/B sky130_fd_sc_hd__xnor2_1
X_6395_ _6795_/CLK _6395_/D vssd1 vssd1 vccd1 vccd1 _6395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5346_ _6625_/Q _5346_/B vssd1 vssd1 vccd1 vccd1 _5347_/A sky130_fd_sc_hd__and2_1
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5277_ _5277_/A vssd1 vssd1 vccd1 vccd1 _6603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4228_ _4228_/A vssd1 vssd1 vccd1 vccd1 _4241_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4159_ _4160_/A _4160_/B _4160_/C vssd1 vssd1 vccd1 vccd1 _4175_/A sky130_fd_sc_hd__o21ai_2
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _3331_/D sky130_fd_sc_hd__clkbuf_4
Xinput45 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
Xinput34 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _3327_/A sky130_fd_sc_hd__clkbuf_2
X_3530_ _3727_/B vssd1 vssd1 vccd1 vccd1 _3755_/B sky130_fd_sc_hd__buf_2
Xinput23 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 _3334_/D sky130_fd_sc_hd__buf_2
Xinput56 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 _4919_/B sky130_fd_sc_hd__clkbuf_4
Xinput67 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_4
X_3461_ _3461_/A vssd1 vssd1 vccd1 vccd1 _6309_/D sky130_fd_sc_hd__clkbuf_1
X_3392_ _3396_/C _3392_/B _3392_/C vssd1 vssd1 vccd1 vccd1 _3393_/A sky130_fd_sc_hd__and3b_1
X_6180_ _6283_/A _6180_/B vssd1 vssd1 vccd1 vccd1 _6180_/X sky130_fd_sc_hd__or2_1
X_5200_ _6701_/Q _6733_/Q _6765_/Q _6797_/Q _5188_/X _5014_/X vssd1 vssd1 vccd1 vccd1
+ _5200_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5131_ _5162_/A vssd1 vssd1 vccd1 vccd1 _5160_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_123_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5062_ _6899_/A _5041_/X _5061_/X _5034_/X vssd1 vssd1 vccd1 vccd1 _6561_/D sky130_fd_sc_hd__o211a_1
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4013_ _4013_/A _4058_/B vssd1 vssd1 vccd1 vccd1 _4017_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5964_ _6248_/A _6286_/A _5964_/C _5964_/D vssd1 vssd1 vccd1 vccd1 _5964_/X sky130_fd_sc_hd__and4b_1
X_4915_ _4915_/A vssd1 vssd1 vccd1 vccd1 _6526_/D sky130_fd_sc_hd__clkbuf_1
X_5895_ _5871_/X _5892_/X _5894_/X _5767_/X vssd1 vssd1 vccd1 vccd1 _5895_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ _4846_/A vssd1 vssd1 vccd1 vccd1 _6485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6516_ _6531_/CLK _6516_/D vssd1 vssd1 vccd1 vccd1 _6516_/Q sky130_fd_sc_hd__dfxtp_1
X_4777_ _4777_/A vssd1 vssd1 vccd1 vccd1 _6454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3728_ _3728_/A _3728_/B vssd1 vssd1 vccd1 vccd1 _3751_/A sky130_fd_sc_hd__or2_1
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3659_ _3659_/A _3755_/C vssd1 vssd1 vccd1 vccd1 _3663_/A sky130_fd_sc_hd__nand2_1
X_6447_ _6789_/CLK _6447_/D vssd1 vssd1 vccd1 vccd1 _6447_/Q sky130_fd_sc_hd__dfxtp_1
X_6378_ _6795_/CLK _6378_/D vssd1 vssd1 vccd1 vccd1 _6378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5329_ _5502_/B _5964_/C _5876_/B vssd1 vssd1 vccd1 vccd1 _5329_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _6364_/Q _4700_/B vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__and2_1
X_5680_ _5735_/A vssd1 vssd1 vccd1 vccd1 _5680_/X sky130_fd_sc_hd__clkbuf_2
X_4631_ _4634_/A _4618_/B _4630_/Y vssd1 vssd1 vccd1 vccd1 _4631_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4562_ _4531_/A _4531_/C _4531_/B vssd1 vssd1 vccd1 vccd1 _4563_/C sky130_fd_sc_hd__a21boi_2
X_4493_ _4493_/A _4493_/B _4493_/C vssd1 vssd1 vccd1 vccd1 _4493_/Y sky130_fd_sc_hd__nand3_2
XFILLER_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6301_ _6509_/CLK _6301_/D vssd1 vssd1 vccd1 vccd1 _6301_/Q sky130_fd_sc_hd__dfxtp_1
X_3513_ _3596_/A _3659_/A _3516_/D _5217_/D vssd1 vssd1 vccd1 vccd1 _3526_/A sky130_fd_sc_hd__nand4_1
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3444_ _3755_/C vssd1 vssd1 vccd1 vccd1 _3810_/B sky130_fd_sc_hd__clkbuf_2
X_6232_ _6800_/Q _6226_/X _6231_/Y _6216_/X vssd1 vssd1 vccd1 vccd1 _6800_/D sky130_fd_sc_hd__o211a_1
X_3375_ _3375_/A _3375_/B vssd1 vssd1 vccd1 vccd1 _6498_/D sky130_fd_sc_hd__nor2_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6775_/Q _6156_/X _6162_/X _6152_/X vssd1 vssd1 vccd1 vccd1 _6775_/D sky130_fd_sc_hd__o211a_1
X_5114_ _6815_/Q _5181_/A vssd1 vssd1 vccd1 vccd1 _5114_/X sky130_fd_sc_hd__or2_1
XFILLER_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6110_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _6095_/A sky130_fd_sc_hd__and2_1
XFILLER_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5011_/X _5043_/X _5044_/X _5019_/X vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__a31o_1
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6996_ _6996_/A _3303_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
XFILLER_92_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5947_ _6107_/A vssd1 vssd1 vccd1 vccd1 _5947_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5878_ _5871_/X _5875_/X _5877_/X vssd1 vssd1 vccd1 vccd1 _5879_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4829_ _4829_/A vssd1 vssd1 vccd1 vccd1 _6477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6886__146 vssd1 vssd1 vccd1 vccd1 _6886__146/HI _6995_/A sky130_fd_sc_hd__conb_1
XFILLER_98_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold1 hold2/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__buf_2
XFILLER_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6781_ _6532_/Q _6781_/D vssd1 vssd1 vccd1 vccd1 _6781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5801_ _6706_/Q _5797_/X _5800_/X _5773_/X vssd1 vssd1 vccd1 vccd1 _6706_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3993_ _4056_/A _4270_/A _3967_/A _3992_/X vssd1 vssd1 vccd1 vccd1 _3994_/A sky130_fd_sc_hd__a31o_1
X_5732_ _6257_/A _5678_/X _5680_/X _5731_/X _5695_/X vssd1 vssd1 vccd1 vccd1 _5732_/X
+ sky130_fd_sc_hd__a221o_1
X_5663_ _5659_/X _5631_/X _5620_/X _5662_/X vssd1 vssd1 vccd1 vccd1 _5663_/X sky130_fd_sc_hd__o211a_1
X_4614_ _4615_/B _4567_/Y _4615_/D _4613_/Y _4590_/B vssd1 vssd1 vccd1 vccd1 _4614_/X
+ sky130_fd_sc_hd__o32a_1
X_5594_ _6453_/Q _5603_/B vssd1 vssd1 vccd1 vccd1 _5594_/X sky130_fd_sc_hd__and2_2
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4545_ _4574_/A _4545_/B _4579_/B _4545_/D vssd1 vssd1 vccd1 vccd1 _4588_/A sky130_fd_sc_hd__and4_1
XFILLER_116_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4476_ _4475_/A _4475_/B _4475_/C vssd1 vssd1 vccd1 vccd1 _4483_/C sky130_fd_sc_hd__a21o_1
X_6215_ _6277_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6215_/X sky130_fd_sc_hd__or2_1
X_3427_ _5214_/D _6504_/Q _3427_/S vssd1 vssd1 vccd1 vccd1 _3428_/A sky130_fd_sc_hd__mux2_1
X_3358_ _3347_/A _3347_/B _6328_/Q vssd1 vssd1 vccd1 vccd1 _3358_/X sky130_fd_sc_hd__o21a_1
X_6146_ _6768_/Q _6142_/X _6145_/X _6051_/X vssd1 vssd1 vccd1 vccd1 _6768_/D sky130_fd_sc_hd__o211a_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3289_ _3292_/A vssd1 vssd1 vccd1 vccd1 _3289_/Y sky130_fd_sc_hd__inv_2
X_6077_ _6754_/Q _6061_/X _6075_/X _6076_/X vssd1 vssd1 vccd1 vccd1 _6078_/B sky130_fd_sc_hd__a22o_1
X_5028_ _6894_/A _4945_/X _5027_/X _4352_/X vssd1 vssd1 vccd1 vccd1 _6556_/D sky130_fd_sc_hd__o211a_1
XFILLER_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6979_ _6979_/A _3283_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4330_ _4576_/C vssd1 vssd1 vccd1 vccd1 _4388_/B sky130_fd_sc_hd__clkbuf_2
X_4261_ _4679_/A vssd1 vssd1 vccd1 vccd1 _4270_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3212_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3212_/Y sky130_fd_sc_hd__inv_2
X_6000_ _6740_/Q _5984_/X _5998_/X _5999_/X vssd1 vssd1 vccd1 vccd1 _6740_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4192_ _4192_/A _4192_/B vssd1 vssd1 vccd1 vccd1 _4198_/B sky130_fd_sc_hd__xnor2_4
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6902_ _6902_/A _3190_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__ebufn_8
XFILLER_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6764_ _6795_/CLK _6764_/D vssd1 vssd1 vccd1 vccd1 _6764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3976_ _4121_/A _4076_/C _4114_/C _4121_/B vssd1 vssd1 vccd1 vccd1 _3977_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5715_ _5560_/X _5698_/X _5699_/X _5714_/X vssd1 vssd1 vccd1 vccd1 _5715_/X sky130_fd_sc_hd__o211a_1
X_6695_ _6809_/CLK _6695_/D vssd1 vssd1 vccd1 vccd1 _6695_/Q sky130_fd_sc_hd__dfxtp_1
X_5646_ _5642_/X _5631_/X _5620_/X _5645_/X vssd1 vssd1 vccd1 vccd1 _5646_/X sky130_fd_sc_hd__o211a_1
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5577_ _6483_/Q vssd1 vssd1 vccd1 vccd1 _6250_/A sky130_fd_sc_hd__buf_2
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4528_ _4540_/A _4540_/B _4540_/C vssd1 vssd1 vccd1 vccd1 _4528_/X sky130_fd_sc_hd__and3_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4459_ _4466_/A _4457_/X _4426_/X _4427_/X vssd1 vssd1 vccd1 vccd1 _4459_/X sky130_fd_sc_hd__o211a_1
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6129_ _6129_/A vssd1 vssd1 vccd1 vccd1 _6764_/D sky130_fd_sc_hd__clkbuf_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3830_ _3827_/X _3828_/X _3825_/Y vssd1 vssd1 vccd1 vccd1 _3831_/B sky130_fd_sc_hd__a21o_1
X_3761_ _3835_/A _3605_/B _3762_/D _3836_/A vssd1 vssd1 vccd1 vccd1 _3763_/A sky130_fd_sc_hd__a22oi_1
X_5500_ _6224_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__nor2_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6480_ _6763_/CLK _6480_/D vssd1 vssd1 vccd1 vccd1 _6480_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3692_ _3692_/A _3692_/B vssd1 vssd1 vccd1 vccd1 _3694_/A sky130_fd_sc_hd__xnor2_2
X_5431_ _5214_/D _3787_/A _5431_/S vssd1 vssd1 vccd1 vccd1 _5432_/B sky130_fd_sc_hd__mux2_1
X_5362_ _5360_/Y _5364_/B _4352_/X vssd1 vssd1 vccd1 vccd1 _6628_/D sky130_fd_sc_hd__o21ai_1
XFILLER_99_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4313_ _6377_/Q vssd1 vssd1 vccd1 vccd1 _4371_/B sky130_fd_sc_hd__clkbuf_2
X_5293_ _5293_/A vssd1 vssd1 vccd1 vccd1 _6610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4244_ _4232_/A _4231_/A _4231_/B _4243_/X vssd1 vssd1 vccd1 vccd1 _4245_/B sky130_fd_sc_hd__a31o_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4175_ _4175_/A vssd1 vssd1 vccd1 vccd1 _4176_/A sky130_fd_sc_hd__inv_2
XFILLER_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6747_ _6532_/Q _6747_/D vssd1 vssd1 vccd1 vccd1 _6747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3959_ _3959_/A _3959_/B vssd1 vssd1 vccd1 vccd1 _4024_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6678_ _6532_/Q _6678_/D vssd1 vssd1 vccd1 vccd1 _6678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5629_ _6682_/Q _5601_/X _5625_/X _5628_/X _5591_/X vssd1 vssd1 vccd1 vccd1 _6682_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_2_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5980_ _6737_/Q _5524_/X _5990_/S vssd1 vssd1 vccd1 vccd1 _5980_/X sky130_fd_sc_hd__mux2_1
X_4931_ _5441_/A vssd1 vssd1 vccd1 vccd1 _4931_/X sky130_fd_sc_hd__buf_4
X_4862_ _6444_/Q _4959_/B vssd1 vssd1 vccd1 vccd1 _4863_/A sky130_fd_sc_hd__and2_1
XFILLER_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6601_ _6667_/CLK _6601_/D vssd1 vssd1 vccd1 vccd1 _6601_/Q sky130_fd_sc_hd__dfxtp_1
X_3813_ _3813_/A _3813_/B _3813_/C vssd1 vssd1 vccd1 vccd1 _3814_/B sky130_fd_sc_hd__nor3_1
XANTENNA_15 _4922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _4566_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4793_ _4793_/A vssd1 vssd1 vccd1 vccd1 _6461_/D sky130_fd_sc_hd__clkbuf_1
X_6532_ _6570_/CLK _6532_/D vssd1 vssd1 vccd1 vccd1 _6532_/Q sky130_fd_sc_hd__dfxtp_4
X_3744_ _3745_/B _3745_/C _3745_/A vssd1 vssd1 vccd1 vccd1 _3778_/C sky130_fd_sc_hd__a21oi_1
XFILLER_20_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3675_ _3592_/X _3631_/B _3629_/X vssd1 vssd1 vccd1 vccd1 _3676_/B sky130_fd_sc_hd__a21oi_2
X_6463_ _6809_/CLK _6463_/D vssd1 vssd1 vccd1 vccd1 _6463_/Q sky130_fd_sc_hd__dfxtp_1
X_5414_ _6604_/Q _6587_/Q _5414_/C _5236_/B vssd1 vssd1 vccd1 vccd1 _5415_/A sky130_fd_sc_hd__or4b_1
XFILLER_114_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6394_ _6795_/CLK _6394_/D vssd1 vssd1 vccd1 vccd1 _6394_/Q sky130_fd_sc_hd__dfxtp_1
X_5345_ _5345_/A vssd1 vssd1 vccd1 vccd1 _6624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5276_ _6603_/Q _5282_/B vssd1 vssd1 vccd1 vccd1 _5277_/A sky130_fd_sc_hd__and2_1
XFILLER_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4227_ _4227_/A vssd1 vssd1 vccd1 vccd1 _4242_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4158_ _4188_/A _4158_/B vssd1 vssd1 vccd1 vccd1 _4160_/C sky130_fd_sc_hd__xnor2_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4089_ _4089_/A _4089_/B _4089_/C vssd1 vssd1 vccd1 vccd1 _4091_/B sky130_fd_sc_hd__nand3_1
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _3331_/C sky130_fd_sc_hd__buf_4
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput35 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _4941_/C sky130_fd_sc_hd__buf_2
Xinput46 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_2
Xinput24 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 _3334_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_116_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput68 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__clkbuf_4
Xinput57 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 _4922_/B sky130_fd_sc_hd__buf_4
XFILLER_115_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3460_ _6309_/Q _6513_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _3461_/A sky130_fd_sc_hd__mux2_1
X_3391_ _6289_/Q _6290_/Q _6291_/Q _6292_/Q vssd1 vssd1 vccd1 vccd1 _3392_/B sky130_fd_sc_hd__a31o_1
X_5130_ _5130_/A vssd1 vssd1 vccd1 vccd1 _6572_/D sky130_fd_sc_hd__clkbuf_1
X_5061_ _5047_/X _5059_/X _5060_/X _5055_/X vssd1 vssd1 vccd1 vccd1 _5061_/X sky130_fd_sc_hd__a31o_1
XFILLER_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4012_ _4183_/B vssd1 vssd1 vccd1 vccd1 _4058_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5963_ _5705_/X _5871_/X _5962_/X vssd1 vssd1 vccd1 vccd1 _5963_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4914_ _4912_/X _6526_/Q _4926_/S vssd1 vssd1 vccd1 vccd1 _4915_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5894_ _6480_/Q _5964_/D _5914_/C vssd1 vssd1 vccd1 vccd1 _5894_/X sky130_fd_sc_hd__and3_1
X_4845_ _6437_/Q _4845_/B vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__and2_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4776_ _6406_/Q _4778_/B vssd1 vssd1 vccd1 vccd1 _4777_/A sky130_fd_sc_hd__and2_1
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6515_ _6531_/CLK _6515_/D vssd1 vssd1 vccd1 vccd1 _6515_/Q sky130_fd_sc_hd__dfxtp_1
X_3727_ _3727_/A _3727_/B _6302_/Q _6301_/Q vssd1 vssd1 vccd1 vccd1 _3728_/B sky130_fd_sc_hd__and4_1
X_3658_ _3679_/B _3679_/C _3679_/A vssd1 vssd1 vccd1 vccd1 _3665_/C sky130_fd_sc_hd__a21o_1
X_6446_ _6789_/CLK _6446_/D vssd1 vssd1 vccd1 vccd1 _6446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6377_ _6795_/CLK _6377_/D vssd1 vssd1 vccd1 vccd1 _6377_/Q sky130_fd_sc_hd__dfxtp_1
X_3589_ _3599_/A _3599_/B vssd1 vssd1 vccd1 vccd1 _3627_/B sky130_fd_sc_hd__xnor2_1
X_5328_ _5880_/A vssd1 vssd1 vccd1 vccd1 _5876_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5259_ _5259_/A vssd1 vssd1 vccd1 vccd1 _6595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _4630_/A _4630_/B vssd1 vssd1 vccd1 vccd1 _4630_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4561_ _4573_/B _4559_/Y _4540_/B _4540_/Y vssd1 vssd1 vccd1 vccd1 _4563_/B sky130_fd_sc_hd__o211a_1
X_6300_ _6504_/CLK _6300_/D vssd1 vssd1 vccd1 vccd1 _6300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4492_ _4493_/B _4493_/C _4493_/A vssd1 vssd1 vccd1 vccd1 _4492_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3512_ _3639_/A _5217_/C _3865_/A _3706_/A vssd1 vssd1 vccd1 vccd1 _3514_/B sky130_fd_sc_hd__a22o_1
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3443_ _6303_/Q vssd1 vssd1 vccd1 vccd1 _3755_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6231_ _6227_/X _6229_/Y _6230_/X vssd1 vssd1 vccd1 vccd1 _6231_/Y sky130_fd_sc_hd__o21ai_1
X_6162_ _6257_/A _6167_/B vssd1 vssd1 vccd1 vccd1 _6162_/X sky130_fd_sc_hd__or2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _6497_/Q _3373_/B _6498_/Q vssd1 vssd1 vccd1 vccd1 _3375_/B sky130_fd_sc_hd__a21oi_1
X_5113_ _5113_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5113_/X sky130_fd_sc_hd__or2_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6757_/Q _6080_/X _6092_/X _6076_/X vssd1 vssd1 vccd1 vccd1 _6094_/B sky130_fd_sc_hd__a22o_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _6804_/Q _5044_/B vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__or2_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6995_ _6995_/A _3302_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
X_5946_ _5946_/A vssd1 vssd1 vccd1 vccd1 _5946_/X sky130_fd_sc_hd__buf_2
XFILLER_53_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5877_ _6720_/Q _5519_/X _5964_/C _5876_/X vssd1 vssd1 vccd1 vccd1 _5877_/X sky130_fd_sc_hd__a22o_1
X_4828_ _6429_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4829_/A sky130_fd_sc_hd__and2_1
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4759_ _6398_/Q _4767_/B vssd1 vssd1 vccd1 vccd1 _4760_/A sky130_fd_sc_hd__and2_1
X_6429_ _6795_/CLK _6429_/D vssd1 vssd1 vccd1 vccd1 _6429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6818__78 vssd1 vssd1 vccd1 vccd1 _6818__78/HI _6927_/A sky130_fd_sc_hd__conb_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6832__92 vssd1 vssd1 vccd1 vccd1 _6832__92/HI _6941_/A sky130_fd_sc_hd__conb_1
X_6780_ _6532_/Q _6780_/D vssd1 vssd1 vccd1 vccd1 _6780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5800_ _6480_/Q _5787_/X _5799_/X _5777_/X _5788_/X vssd1 vssd1 vccd1 vccd1 _5800_/X
+ sky130_fd_sc_hd__a221o_1
X_3992_ _3992_/A _4268_/A _3992_/C vssd1 vssd1 vccd1 vccd1 _3992_/X sky130_fd_sc_hd__and3_1
XFILLER_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5731_ _5593_/X _5729_/X _5757_/S vssd1 vssd1 vccd1 vccd1 _5731_/X sky130_fd_sc_hd__mux2_1
X_5662_ _5670_/A _5662_/B vssd1 vssd1 vccd1 vccd1 _5662_/X sky130_fd_sc_hd__or2_1
XFILLER_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4613_ _4613_/A _4613_/B vssd1 vssd1 vccd1 vccd1 _4613_/Y sky130_fd_sc_hd__nor2_1
X_5593_ _6469_/Q vssd1 vssd1 vccd1 vccd1 _5593_/X sky130_fd_sc_hd__clkbuf_4
X_4544_ _4574_/A _4579_/B _4545_/D _4545_/B vssd1 vssd1 vccd1 vccd1 _4546_/A sky130_fd_sc_hd__a22oi_1
XFILLER_89_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6214_ _6795_/Q _6207_/X _6213_/X _6203_/X vssd1 vssd1 vccd1 vccd1 _6795_/D sky130_fd_sc_hd__o211a_1
X_4475_ _4475_/A _4475_/B _4475_/C vssd1 vssd1 vccd1 vccd1 _4483_/B sky130_fd_sc_hd__nand3_1
XFILLER_116_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3426_ _3722_/B vssd1 vssd1 vccd1 vccd1 _5214_/D sky130_fd_sc_hd__buf_2
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3357_ _6011_/A vssd1 vssd1 vccd1 vccd1 _3357_/X sky130_fd_sc_hd__clkbuf_4
X_6145_ _6229_/A _6154_/B vssd1 vssd1 vccd1 vccd1 _6145_/X sky130_fd_sc_hd__or2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6076_ _6102_/A vssd1 vssd1 vccd1 vccd1 _6076_/X sky130_fd_sc_hd__clkbuf_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3288_ _3292_/A vssd1 vssd1 vccd1 vccd1 _3288_/Y sky130_fd_sc_hd__inv_2
X_5027_ _5011_/X _5023_/X _5026_/X _5019_/X vssd1 vssd1 vccd1 vccd1 _5027_/X sky130_fd_sc_hd__a31o_1
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6978_ _6978_/A _3282_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5929_ _6728_/Q _5918_/X _5928_/X _5904_/X vssd1 vssd1 vccd1 vccd1 _6728_/D sky130_fd_sc_hd__o211a_1
XFILLER_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6853__113 vssd1 vssd1 vccd1 vccd1 _6853__113/HI _6962_/A sky130_fd_sc_hd__conb_1
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4260_ _5458_/A vssd1 vssd1 vccd1 vccd1 _4679_/A sky130_fd_sc_hd__buf_4
X_3211_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3211_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4191_ _4212_/A _4212_/B vssd1 vssd1 vccd1 vccd1 _4192_/B sky130_fd_sc_hd__xor2_4
XFILLER_94_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6901_ _6901_/A _3189_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__ebufn_8
XFILLER_63_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6763_ _6763_/CLK _6763_/D vssd1 vssd1 vccd1 vccd1 _6763_/Q sky130_fd_sc_hd__dfxtp_1
X_3975_ _6352_/Q vssd1 vssd1 vccd1 vccd1 _4114_/C sky130_fd_sc_hd__clkbuf_2
X_5714_ _5765_/A _5714_/B vssd1 vssd1 vccd1 vccd1 _5714_/X sky130_fd_sc_hd__or2_1
X_6694_ _6809_/CLK _6694_/D vssd1 vssd1 vccd1 vccd1 _6694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5645_ _5670_/A _5645_/B vssd1 vssd1 vccd1 vccd1 _5645_/X sky130_fd_sc_hd__or2_1
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5576_ _5570_/X _5525_/X _5571_/X _5575_/X vssd1 vssd1 vccd1 vccd1 _5576_/X sky130_fd_sc_hd__o211a_1
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4527_ _4540_/B _4540_/C _4540_/A vssd1 vssd1 vccd1 vccd1 _4527_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4458_ _4426_/X _4427_/X _4466_/A _4457_/X vssd1 vssd1 vccd1 vccd1 _4458_/Y sky130_fd_sc_hd__a211oi_2
X_3409_ _3409_/A vssd1 vssd1 vccd1 vccd1 _6296_/D sky130_fd_sc_hd__clkbuf_1
X_4389_ _4283_/A _4595_/C _4363_/A _4388_/X vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__a31o_1
XFILLER_86_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6128_ _6132_/A _6128_/B vssd1 vssd1 vccd1 vccd1 _6129_/A sky130_fd_sc_hd__and2_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6059_ _6059_/A _6068_/A vssd1 vssd1 vccd1 vccd1 _6059_/X sky130_fd_sc_hd__or2_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3760_ _6655_/Q vssd1 vssd1 vccd1 vccd1 _3836_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3691_ _3691_/A _3691_/B vssd1 vssd1 vccd1 vccd1 _3692_/B sky130_fd_sc_hd__nor2_1
X_5430_ _5430_/A vssd1 vssd1 vccd1 vccd1 _6651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5361_ _5882_/A _6224_/B _5971_/B vssd1 vssd1 vccd1 vccd1 _5364_/B sky130_fd_sc_hd__and3_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5292_ _6610_/Q _5294_/B vssd1 vssd1 vccd1 vccd1 _5293_/A sky130_fd_sc_hd__and2_1
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4312_ _4354_/C _4312_/B vssd1 vssd1 vccd1 vccd1 _4319_/A sky130_fd_sc_hd__or2_1
XFILLER_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4243_ _4243_/A _4247_/B vssd1 vssd1 vccd1 vccd1 _4243_/X sky130_fd_sc_hd__and2_1
XFILLER_113_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _4195_/B _4174_/B vssd1 vssd1 vccd1 vccd1 _6368_/D sky130_fd_sc_hd__nor2_1
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6815_ _6532_/Q _6815_/D vssd1 vssd1 vccd1 vccd1 _6815_/Q sky130_fd_sc_hd__dfxtp_1
X_6746_ _6532_/Q _6746_/D vssd1 vssd1 vccd1 vccd1 _6746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3958_ _4056_/A _4268_/A _3940_/A _3957_/X vssd1 vssd1 vccd1 vccd1 _3985_/A sky130_fd_sc_hd__a31o_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6677_ _6809_/CLK _6677_/D vssd1 vssd1 vccd1 vccd1 _6677_/Q sky130_fd_sc_hd__dfxtp_1
X_3889_ _3889_/A _4257_/A _5008_/B vssd1 vssd1 vccd1 vccd1 _3890_/A sky130_fd_sc_hd__and3_1
X_5628_ _6270_/A _5589_/X _5627_/X _5616_/X vssd1 vssd1 vccd1 vccd1 _5628_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5559_ _6675_/Q _5551_/X _5556_/X _5558_/X _5540_/X vssd1 vssd1 vccd1 vccd1 _6675_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_120_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4930_ _4930_/A vssd1 vssd1 vccd1 vccd1 _6531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4861_ _4861_/A vssd1 vssd1 vccd1 vccd1 _6491_/D sky130_fd_sc_hd__clkbuf_1
X_6600_ _6667_/CLK _6600_/D vssd1 vssd1 vccd1 vccd1 _6600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3812_ _3813_/A _3813_/B _3813_/C vssd1 vssd1 vccd1 vccd1 _3851_/A sky130_fd_sc_hd__o21a_1
XANTENNA_16 _4928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4792_ _6413_/Q _4800_/B vssd1 vssd1 vccd1 vccd1 _4793_/A sky130_fd_sc_hd__and2_1
XANTENNA_27 _5570_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6531_ _6531_/CLK _6531_/D vssd1 vssd1 vccd1 vccd1 _6531_/Q sky130_fd_sc_hd__dfxtp_1
X_3743_ _3709_/A _3709_/C _3709_/B vssd1 vssd1 vccd1 vccd1 _3745_/A sky130_fd_sc_hd__a21bo_1
X_3674_ _3674_/A _3673_/X vssd1 vssd1 vccd1 vccd1 _3676_/A sky130_fd_sc_hd__or2b_1
X_6462_ _6809_/CLK _6462_/D vssd1 vssd1 vccd1 vccd1 _6462_/Q sky130_fd_sc_hd__dfxtp_2
X_5413_ _5413_/A vssd1 vssd1 vccd1 vccd1 _6647_/D sky130_fd_sc_hd__clkbuf_1
X_6393_ _6795_/CLK _6393_/D vssd1 vssd1 vccd1 vccd1 _6393_/Q sky130_fd_sc_hd__dfxtp_1
X_5344_ _6624_/Q _5346_/B vssd1 vssd1 vccd1 vccd1 _5345_/A sky130_fd_sc_hd__and2_1
XFILLER_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5275_ _5275_/A vssd1 vssd1 vccd1 vccd1 _6602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4226_ _4203_/A _4203_/B _4201_/B vssd1 vssd1 vccd1 vccd1 _4232_/A sky130_fd_sc_hd__o21ai_2
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4157_ _4157_/A _4189_/A vssd1 vssd1 vccd1 vccd1 _4158_/B sky130_fd_sc_hd__xnor2_2
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4088_ _4089_/B _4089_/C _4089_/A vssd1 vssd1 vccd1 vccd1 _4091_/A sky130_fd_sc_hd__a21o_1
XFILLER_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6729_ _6799_/CLK _6729_/D vssd1 vssd1 vccd1 vccd1 _6729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput36 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_4
Xinput14 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _3326_/A sky130_fd_sc_hd__clkbuf_2
Xinput25 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _3326_/D sky130_fd_sc_hd__buf_2
Xinput69 wbs_we_i vssd1 vssd1 vccd1 vccd1 _3324_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
Xinput58 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_2
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3390_ _6292_/Q _6291_/Q _3390_/C vssd1 vssd1 vccd1 vccd1 _3396_/C sky130_fd_sc_hd__and3_1
XFILLER_96_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5060_ _6806_/Q _5078_/B vssd1 vssd1 vccd1 vccd1 _5060_/X sky130_fd_sc_hd__or2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4011_ _6356_/Q vssd1 vssd1 vccd1 vccd1 _4183_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ _6735_/Q _5667_/X _5962_/S vssd1 vssd1 vccd1 vccd1 _5962_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4913_ _4929_/S vssd1 vssd1 vccd1 vccd1 _4926_/S sky130_fd_sc_hd__buf_2
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5893_ _5922_/A vssd1 vssd1 vccd1 vccd1 _5914_/C sky130_fd_sc_hd__clkbuf_1
X_4844_ _4844_/A vssd1 vssd1 vccd1 vccd1 _6484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4775_ _4775_/A vssd1 vssd1 vccd1 vccd1 _6453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6514_ _6522_/CLK _6514_/D vssd1 vssd1 vccd1 vccd1 _6514_/Q sky130_fd_sc_hd__dfxtp_1
X_3726_ _3690_/B _3755_/D _3789_/C _3753_/A vssd1 vssd1 vccd1 vccd1 _3728_/A sky130_fd_sc_hd__a22oi_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6445_ _6795_/CLK _6445_/D vssd1 vssd1 vccd1 vccd1 _6445_/Q sky130_fd_sc_hd__dfxtp_1
X_3657_ _3679_/A _3679_/B _3679_/C vssd1 vssd1 vccd1 vccd1 _3665_/B sky130_fd_sc_hd__nand3_1
X_6376_ _6795_/CLK _6376_/D vssd1 vssd1 vccd1 vccd1 _6376_/Q sky130_fd_sc_hd__dfxtp_1
X_3588_ _3614_/A _3588_/B vssd1 vssd1 vccd1 vccd1 _3599_/B sky130_fd_sc_hd__nor2_2
X_5327_ _6621_/Q vssd1 vssd1 vccd1 vccd1 _5880_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5258_ _6595_/Q _5260_/B vssd1 vssd1 vccd1 vccd1 _5259_/A sky130_fd_sc_hd__and2_1
XFILLER_102_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5189_ _6699_/Q _6731_/Q _6763_/Q _6795_/Q _5188_/X _5169_/X vssd1 vssd1 vccd1 vccd1
+ _5189_/X sky130_fd_sc_hd__mux4_1
X_4209_ _4210_/A _4210_/B vssd1 vssd1 vccd1 vccd1 _4211_/A sky130_fd_sc_hd__and2_1
XFILLER_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4560_ _4540_/B _4540_/Y _4573_/B _4559_/Y vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__a211oi_4
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4491_ _4531_/A _4491_/B vssd1 vssd1 vccd1 vccd1 _4493_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3511_ _3596_/A vssd1 vssd1 vccd1 vccd1 _3706_/A sky130_fd_sc_hd__clkbuf_2
X_6230_ _6264_/A vssd1 vssd1 vccd1 vccd1 _6230_/X sky130_fd_sc_hd__buf_2
X_3442_ _3442_/A vssd1 vssd1 vccd1 vccd1 _6302_/D sky130_fd_sc_hd__clkbuf_1
X_3373_ _6497_/Q _3373_/B vssd1 vssd1 vccd1 vccd1 _6497_/D sky130_fd_sc_hd__xor2_1
X_6161_ _6774_/Q _6156_/X _6160_/X _6152_/X vssd1 vssd1 vccd1 vccd1 _6774_/D sky130_fd_sc_hd__o211a_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _6687_/Q _6719_/Q _6751_/Q _6783_/Q _5188_/A _4949_/A vssd1 vssd1 vccd1 vccd1
+ _5113_/B sky130_fd_sc_hd__mux4_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6467_/Q _6081_/X _6070_/X _6087_/X _6483_/Q vssd1 vssd1 vccd1 vccd1 _6092_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5043_/A _5043_/B vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__or2_1
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6994_ _6994_/A _3301_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5945_ _6731_/Q _5918_/X _5944_/X _5933_/X vssd1 vssd1 vccd1 vccd1 _6731_/D sky130_fd_sc_hd__o211a_1
X_5876_ _6268_/A _5876_/B _6478_/Q _5880_/B vssd1 vssd1 vccd1 vccd1 _5876_/X sky130_fd_sc_hd__and4b_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4827_ _4827_/A vssd1 vssd1 vccd1 vccd1 _6476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4758_ _4791_/A vssd1 vssd1 vccd1 vccd1 _4767_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3709_ _3709_/A _3709_/B _3709_/C vssd1 vssd1 vccd1 vccd1 _3709_/X sky130_fd_sc_hd__and3_1
X_4689_ _4689_/A vssd1 vssd1 vccd1 vccd1 _6415_/D sky130_fd_sc_hd__clkbuf_1
X_6428_ _6763_/CLK _6428_/D vssd1 vssd1 vccd1 vccd1 _6428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6359_ _6763_/CLK _6359_/D vssd1 vssd1 vccd1 vccd1 _6359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3991_ _4151_/B vssd1 vssd1 vccd1 vccd1 _4270_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5730_ _5771_/S vssd1 vssd1 vccd1 vccd1 _5757_/S sky130_fd_sc_hd__buf_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5661_ _6686_/Q _5660_/X _5661_/S vssd1 vssd1 vccd1 vccd1 _5662_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4612_ _4634_/A _4612_/B vssd1 vssd1 vccd1 vccd1 _4612_/Y sky130_fd_sc_hd__nand2_1
X_5592_ _6678_/Q _5551_/X _5587_/X _5590_/X _5591_/X vssd1 vssd1 vccd1 vccd1 _6678_/D
+ sky130_fd_sc_hd__o221a_1
X_4543_ _4543_/A vssd1 vssd1 vccd1 vccd1 _4574_/A sky130_fd_sc_hd__clkbuf_2
X_4474_ _4436_/A _4436_/B _4436_/C vssd1 vssd1 vccd1 vccd1 _4475_/C sky130_fd_sc_hd__a21bo_1
X_6213_ _6273_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6213_/X sky130_fd_sc_hd__or2_1
X_3425_ _3789_/D vssd1 vssd1 vccd1 vccd1 _3722_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_112_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3356_ _5406_/C vssd1 vssd1 vccd1 vccd1 _6011_/A sky130_fd_sc_hd__buf_2
X_6144_ _6182_/B vssd1 vssd1 vccd1 vccd1 _6154_/B sky130_fd_sc_hd__clkbuf_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3305_/A vssd1 vssd1 vccd1 vccd1 _3292_/A sky130_fd_sc_hd__buf_12
XFILLER_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6464_/Q _5947_/X _6070_/X _6138_/S _6480_/Q vssd1 vssd1 vccd1 vccd1 _6075_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5026_ _6801_/Q _5044_/B vssd1 vssd1 vccd1 vccd1 _5026_/X sky130_fd_sc_hd__or2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6977_ _6977_/A _3280_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5928_ _5906_/X _5926_/X _5927_/X _5915_/X vssd1 vssd1 vccd1 vccd1 _5928_/X sky130_fd_sc_hd__a211o_1
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5859_ _6718_/Q _5660_/X _5859_/S vssd1 vssd1 vccd1 vccd1 _5859_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3210_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3210_/Y sky130_fd_sc_hd__inv_2
X_4190_ _4188_/Y _4158_/B _4189_/X vssd1 vssd1 vccd1 vccd1 _4212_/B sky130_fd_sc_hd__a21bo_1
XFILLER_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6900_ _6900_/A _3187_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__ebufn_8
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6762_ _6763_/CLK _6762_/D vssd1 vssd1 vccd1 vccd1 _6762_/Q sky130_fd_sc_hd__dfxtp_1
X_3974_ _6353_/Q vssd1 vssd1 vccd1 vccd1 _3998_/D sky130_fd_sc_hd__clkbuf_2
X_6693_ _6809_/CLK _6693_/D vssd1 vssd1 vccd1 vccd1 _6693_/Q sky130_fd_sc_hd__dfxtp_1
X_5713_ _6692_/Q _5561_/X _5724_/S vssd1 vssd1 vccd1 vccd1 _5714_/B sky130_fd_sc_hd__mux2_1
X_5644_ _6684_/Q _5643_/X _5661_/S vssd1 vssd1 vccd1 vccd1 _5645_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6509_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_5575_ _5575_/A _5575_/B vssd1 vssd1 vccd1 vccd1 _5575_/X sky130_fd_sc_hd__or2_1
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4526_ _4333_/A _4595_/D _4481_/B _4480_/B vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__a31o_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4457_ _4454_/Y _4455_/X _4428_/B _4428_/Y vssd1 vssd1 vccd1 vccd1 _4457_/X sky130_fd_sc_hd__o211a_1
X_3408_ _3865_/A _6500_/Q _3427_/S vssd1 vssd1 vccd1 vccd1 _3409_/A sky130_fd_sc_hd__mux2_1
X_4388_ _4499_/A _4388_/B _4388_/C vssd1 vssd1 vccd1 vccd1 _4388_/X sky130_fd_sc_hd__and3_1
X_6127_ _6764_/Q _6106_/X _6126_/X _5406_/C vssd1 vssd1 vccd1 vccd1 _6128_/B sky130_fd_sc_hd__a22o_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _5441_/A vssd1 vssd1 vccd1 vccd1 _5422_/A sky130_fd_sc_hd__buf_4
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6058_ _6058_/A _6062_/C vssd1 vssd1 vccd1 vccd1 _6058_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5009_ _5009_/A vssd1 vssd1 vccd1 vccd1 _6553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6876__136 vssd1 vssd1 vccd1 vccd1 _6876__136/HI _6985_/A sky130_fd_sc_hd__conb_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3690_ _3727_/A _3690_/B _3789_/C _3789_/D vssd1 vssd1 vccd1 vccd1 _3691_/B sky130_fd_sc_hd__and4_1
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5360_ _5797_/A _5971_/B _5873_/A vssd1 vssd1 vccd1 vccd1 _5360_/Y sky130_fd_sc_hd__a21oi_1
X_5291_ _5291_/A vssd1 vssd1 vccd1 vccd1 _6609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4311_ _4545_/B _4373_/D _4296_/C _4477_/A vssd1 vssd1 vccd1 vccd1 _4312_/B sky130_fd_sc_hd__a22oi_1
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4242_ _4242_/A _4275_/A _4242_/C vssd1 vssd1 vccd1 vccd1 _4245_/A sky130_fd_sc_hd__and3_1
X_4173_ _4220_/B _4172_/B _5001_/A vssd1 vssd1 vccd1 vccd1 _4174_/B sky130_fd_sc_hd__a21o_1
XFILLER_95_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6814_ _6532_/Q _6814_/D vssd1 vssd1 vccd1 vccd1 _6814_/Q sky130_fd_sc_hd__dfxtp_1
X_6745_ _6532_/Q _6745_/D vssd1 vssd1 vccd1 vccd1 _6745_/Q sky130_fd_sc_hd__dfxtp_1
X_3957_ _4103_/A _4266_/A _3957_/C vssd1 vssd1 vccd1 vccd1 _3957_/X sky130_fd_sc_hd__and3_1
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6676_ _6809_/CLK _6676_/D vssd1 vssd1 vccd1 vccd1 _6676_/Q sky130_fd_sc_hd__dfxtp_1
X_3888_ _3979_/D vssd1 vssd1 vccd1 vccd1 _4257_/A sky130_fd_sc_hd__clkbuf_2
X_5627_ _6269_/A vssd1 vssd1 vccd1 vccd1 _5627_/X sky130_fd_sc_hd__clkbuf_2
X_5558_ _6240_/A _5534_/X _6286_/B _5538_/X vssd1 vssd1 vccd1 vccd1 _5558_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4509_ _6671_/Q _6376_/Q _6377_/Q _4510_/B vssd1 vssd1 vccd1 vccd1 _4512_/C sky130_fd_sc_hd__a22o_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5489_ _6317_/Q _4597_/A _5496_/S vssd1 vssd1 vccd1 vccd1 _5490_/B sky130_fd_sc_hd__mux2_1
XFILLER_120_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4860_ _6443_/Q _4959_/B vssd1 vssd1 vccd1 vccd1 _4861_/A sky130_fd_sc_hd__and2_1
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3811_ _3811_/A _3811_/B vssd1 vssd1 vccd1 vccd1 _3813_/C sky130_fd_sc_hd__xor2_1
XFILLER_33_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6530_ _6554_/CLK _6530_/D vssd1 vssd1 vccd1 vccd1 _6530_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_28 _6492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4791_ _4791_/A vssd1 vssd1 vccd1 vccd1 _4800_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3742_ _3741_/B _3741_/C _3741_/A vssd1 vssd1 vccd1 vccd1 _3745_/C sky130_fd_sc_hd__a21o_1
X_3673_ _3671_/X _3629_/A _3669_/X _3670_/Y vssd1 vssd1 vccd1 vccd1 _3673_/X sky130_fd_sc_hd__a211o_1
X_6461_ _6789_/CLK _6461_/D vssd1 vssd1 vccd1 vccd1 _6461_/Q sky130_fd_sc_hd__dfxtp_1
X_5412_ _6647_/Q _5412_/B vssd1 vssd1 vccd1 vccd1 _5413_/A sky130_fd_sc_hd__and2_1
X_6392_ _6795_/CLK _6392_/D vssd1 vssd1 vccd1 vccd1 _6392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5343_ _6224_/A _5342_/X _5331_/X vssd1 vssd1 vccd1 vccd1 _6623_/D sky130_fd_sc_hd__o21a_1
X_5274_ _6602_/Q _5282_/B vssd1 vssd1 vccd1 vccd1 _5275_/A sky130_fd_sc_hd__and2_1
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4225_ _4214_/B _4225_/B vssd1 vssd1 vccd1 vccd1 _4235_/A sky130_fd_sc_hd__and2b_1
XFILLER_101_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4156_ _4156_/A _4156_/B vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__and2_1
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _4087_/A _4087_/B vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__xnor2_2
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4989_ _6545_/Q _4986_/B _6546_/Q vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__a21oi_1
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6728_ _6799_/CLK _6728_/D vssd1 vssd1 vccd1 vccd1 _6728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6659_ _6795_/CLK _6659_/D vssd1 vssd1 vccd1 vccd1 _6659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput37 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_2
Xinput26 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_2
Xinput15 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _3330_/B sky130_fd_sc_hd__buf_2
XFILLER_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput59 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 _4925_/B sky130_fd_sc_hd__buf_6
Xinput48 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6839__99 vssd1 vssd1 vccd1 vccd1 _6839__99/HI _6948_/A sky130_fd_sc_hd__conb_1
XFILLER_96_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4010_ _4009_/B _4009_/C _4009_/A vssd1 vssd1 vccd1 vccd1 _4019_/C sky130_fd_sc_hd__a21o_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5961_ _6003_/A _5961_/B vssd1 vssd1 vccd1 vccd1 _5962_/S sky130_fd_sc_hd__nor2_1
XFILLER_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ _4919_/A _4912_/B vssd1 vssd1 vccd1 vccd1 _4912_/X sky130_fd_sc_hd__and2_1
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5892_ _5542_/X _5889_/X _5891_/X _5874_/X _6722_/Q vssd1 vssd1 vccd1 vccd1 _5892_/X
+ sky130_fd_sc_hd__a32o_1
X_4843_ _6436_/Q _4845_/B vssd1 vssd1 vccd1 vccd1 _4844_/A sky130_fd_sc_hd__and2_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4774_ _6405_/Q _4778_/B vssd1 vssd1 vccd1 vccd1 _4775_/A sky130_fd_sc_hd__and2_1
X_6513_ _6522_/CLK _6513_/D vssd1 vssd1 vccd1 vccd1 _6513_/Q sky130_fd_sc_hd__dfxtp_1
X_3725_ _3724_/A _3765_/B _3724_/C vssd1 vssd1 vccd1 vccd1 _3752_/B sky130_fd_sc_hd__a21oi_1
XFILLER_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6444_ _6795_/CLK _6444_/D vssd1 vssd1 vccd1 vccd1 _6444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3656_ _3656_/A _3656_/B _3656_/C vssd1 vssd1 vccd1 vccd1 _3679_/C sky130_fd_sc_hd__nand3_1
X_6375_ _6795_/CLK _6375_/D vssd1 vssd1 vccd1 vccd1 _6375_/Q sky130_fd_sc_hd__dfxtp_1
X_3587_ _3586_/B _3586_/C _3586_/A vssd1 vssd1 vccd1 vccd1 _3588_/B sky130_fd_sc_hd__o21a_1
X_5326_ _5502_/B _5964_/C _5325_/Y vssd1 vssd1 vccd1 vccd1 _6620_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5257_ _5257_/A vssd1 vssd1 vccd1 vccd1 _6594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4208_ _4177_/A _4275_/A _4187_/B _4207_/X vssd1 vssd1 vccd1 vccd1 _4210_/B sky130_fd_sc_hd__a31oi_2
X_5188_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__buf_2
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4139_ _4169_/A _4169_/B _4169_/C vssd1 vssd1 vccd1 vccd1 _4140_/B sky130_fd_sc_hd__nand3_1
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3510_ _3661_/A vssd1 vssd1 vccd1 vccd1 _3596_/A sky130_fd_sc_hd__clkbuf_2
X_4490_ _4296_/A _4597_/B _4442_/B _4487_/Y vssd1 vssd1 vccd1 vccd1 _4491_/B sky130_fd_sc_hd__a211oi_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3441_ _3879_/A _6506_/Q _3451_/S vssd1 vssd1 vccd1 vccd1 _3442_/A sky130_fd_sc_hd__mux2_1
X_3372_ _3373_/B _3372_/B vssd1 vssd1 vccd1 vccd1 _6496_/D sky130_fd_sc_hd__nor2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6160_ _6253_/A _6167_/B vssd1 vssd1 vccd1 vccd1 _6160_/X sky130_fd_sc_hd__or2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5111_ _6907_/A _5041_/A _5110_/X _5100_/X vssd1 vssd1 vccd1 vccd1 _6569_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6091_/A vssd1 vssd1 vccd1 vccd1 _6756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _6676_/Q _6708_/Q _6740_/Q _6772_/Q _5012_/X _5029_/X vssd1 vssd1 vccd1 vccd1
+ _5043_/B sky130_fd_sc_hd__mux4_1
XFILLER_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6993_ _6993_/A _3300_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5944_ _5935_/X _5942_/X _5943_/X _5687_/X vssd1 vssd1 vccd1 vccd1 _5944_/X sky130_fd_sc_hd__a211o_1
X_5875_ _5506_/X _5364_/X _5874_/X _6720_/Q vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4826_ _6428_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4827_/A sky130_fd_sc_hd__and2_1
X_4757_ _4757_/A vssd1 vssd1 vccd1 vccd1 _6445_/D sky130_fd_sc_hd__clkbuf_1
X_3708_ _3709_/B _3709_/C _3709_/A vssd1 vssd1 vccd1 vccd1 _3708_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4688_ _6359_/Q _4688_/B vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__and2_1
X_6427_ _6763_/CLK _6427_/D vssd1 vssd1 vccd1 vccd1 _6427_/Q sky130_fd_sc_hd__dfxtp_1
X_3639_ _3639_/A _5214_/B _3639_/C vssd1 vssd1 vccd1 vccd1 _3639_/X sky130_fd_sc_hd__and3_1
X_6358_ _6763_/CLK _6358_/D vssd1 vssd1 vccd1 vccd1 _6358_/Q sky130_fd_sc_hd__dfxtp_1
X_5309_ _5309_/A vssd1 vssd1 vccd1 vccd1 _6617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6289_ _6584_/CLK _6289_/D vssd1 vssd1 vccd1 vccd1 _6289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3990_ _3990_/A vssd1 vssd1 vccd1 vccd1 _6363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5660_ _6460_/Q _5660_/B vssd1 vssd1 vccd1 vccd1 _5660_/X sky130_fd_sc_hd__and2_2
XFILLER_90_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4611_ _4611_/A _4611_/B vssd1 vssd1 vccd1 vccd1 _4612_/B sky130_fd_sc_hd__nand2_1
X_5591_ _5707_/A vssd1 vssd1 vccd1 vccd1 _5591_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4542_ _4557_/A _4542_/B _4520_/X vssd1 vssd1 vccd1 vccd1 _4557_/B sky130_fd_sc_hd__nor3b_1
X_4473_ _4473_/A _4473_/B _4473_/C vssd1 vssd1 vccd1 vccd1 _4475_/B sky130_fd_sc_hd__nand3_1
X_6212_ _6794_/Q _6207_/X _6211_/X _6203_/X vssd1 vssd1 vccd1 vccd1 _6794_/D sky130_fd_sc_hd__o211a_1
X_3424_ _6300_/Q vssd1 vssd1 vccd1 vccd1 _3789_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6143_ _6143_/A _6143_/B vssd1 vssd1 vccd1 vccd1 _6182_/B sky130_fd_sc_hd__or2_4
X_3355_ _6102_/A vssd1 vssd1 vccd1 vccd1 _5406_/C sky130_fd_sc_hd__clkbuf_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6074_ _6074_/A vssd1 vssd1 vccd1 vccd1 _6753_/D sky130_fd_sc_hd__clkbuf_1
X_3286_ _3286_/A vssd1 vssd1 vccd1 vccd1 _3286_/Y sky130_fd_sc_hd__inv_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5025_ _5086_/A vssd1 vssd1 vccd1 vccd1 _5044_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6823__83 vssd1 vssd1 vccd1 vccd1 _6823__83/HI _6932_/A sky130_fd_sc_hd__conb_1
XFILLER_81_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6976_ _6976_/A _3279_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5927_ _6486_/Q _5931_/B _5943_/C vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__and3_1
X_5858_ _6717_/Q _5850_/X _5857_/X _5838_/X vssd1 vssd1 vccd1 vccd1 _6717_/D sky130_fd_sc_hd__o211a_1
X_5789_ _5777_/X _5784_/X _5787_/X _6229_/A _5788_/X vssd1 vssd1 vccd1 vccd1 _5789_/X
+ sky130_fd_sc_hd__a221o_1
X_4809_ _4809_/A vssd1 vssd1 vccd1 vccd1 _6468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6761_ _6763_/CLK _6761_/D vssd1 vssd1 vccd1 vccd1 _6761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5712_ _6691_/Q _3357_/X _5711_/X _5690_/X vssd1 vssd1 vccd1 vccd1 _6691_/D sky130_fd_sc_hd__o211a_1
X_3973_ _4123_/A _4266_/A _3970_/Y _3972_/X vssd1 vssd1 vccd1 vccd1 _3973_/X sky130_fd_sc_hd__o2bb2a_1
X_6692_ _6789_/CLK _6692_/D vssd1 vssd1 vccd1 vccd1 _6692_/Q sky130_fd_sc_hd__dfxtp_1
X_5643_ _6458_/Q _5652_/B vssd1 vssd1 vccd1 vccd1 _5643_/X sky130_fd_sc_hd__and2_2
XFILLER_31_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5574_ _6677_/Q _5572_/X _5612_/S vssd1 vssd1 vccd1 vccd1 _5575_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4525_ _4524_/A _4524_/B _4524_/C vssd1 vssd1 vccd1 vccd1 _4540_/C sky130_fd_sc_hd__a21o_1
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4456_ _4428_/B _4428_/Y _4454_/Y _4455_/X vssd1 vssd1 vccd1 vccd1 _4466_/A sky130_fd_sc_hd__a211oi_4
X_4387_ _5162_/A vssd1 vssd1 vccd1 vccd1 _5129_/A sky130_fd_sc_hd__buf_2
X_3407_ _3499_/S vssd1 vssd1 vccd1 vccd1 _3427_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_49_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3338_ _5284_/A vssd1 vssd1 vccd1 vccd1 _5441_/A sky130_fd_sc_hd__clkbuf_4
X_6126_ _6474_/Q _6107_/X _6070_/A _6113_/X _6490_/Q vssd1 vssd1 vccd1 vccd1 _6126_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _3281_/A vssd1 vssd1 vccd1 vccd1 _3274_/A sky130_fd_sc_hd__buf_12
X_6057_ _6751_/Q _5380_/X _6055_/X _6056_/X _4931_/X vssd1 vssd1 vccd1 vccd1 _6751_/D
+ sky130_fd_sc_hd__o221a_1
X_5008_ _5008_/A _5008_/B _5008_/C vssd1 vssd1 vccd1 vccd1 _5009_/A sky130_fd_sc_hd__and3_1
XFILLER_54_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6959_ _6959_/A _3260_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5290_ _6609_/Q _5294_/B vssd1 vssd1 vccd1 vccd1 _5291_/A sky130_fd_sc_hd__and2_1
XFILLER_99_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4310_ _4517_/B vssd1 vssd1 vccd1 vccd1 _4545_/B sky130_fd_sc_hd__buf_2
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4241_ _4241_/A _4273_/A vssd1 vssd1 vccd1 vccd1 _4242_/C sky130_fd_sc_hd__nand2_1
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4172_ _4220_/B _4172_/B vssd1 vssd1 vccd1 vccd1 _4195_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6813_ _6532_/Q _6813_/D vssd1 vssd1 vccd1 vccd1 _6813_/Q sky130_fd_sc_hd__dfxtp_1
X_6744_ _6532_/Q _6744_/D vssd1 vssd1 vccd1 vccd1 _6744_/Q sky130_fd_sc_hd__dfxtp_1
X_3956_ _3956_/A vssd1 vssd1 vccd1 vccd1 _3988_/A sky130_fd_sc_hd__inv_2
X_6675_ _6809_/CLK _6675_/D vssd1 vssd1 vccd1 vccd1 _6675_/Q sky130_fd_sc_hd__dfxtp_1
X_5626_ _6488_/Q vssd1 vssd1 vccd1 vccd1 _6270_/A sky130_fd_sc_hd__buf_4
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3887_ _4039_/C vssd1 vssd1 vccd1 vccd1 _3979_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5557_ _6481_/Q vssd1 vssd1 vccd1 vccd1 _6240_/A sky130_fd_sc_hd__buf_2
XFILLER_117_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4508_ _4505_/X _4615_/A _4507_/Y vssd1 vssd1 vccd1 vccd1 _6390_/D sky130_fd_sc_hd__o21a_1
X_5488_ _5488_/A vssd1 vssd1 vccd1 vccd1 _6668_/D sky130_fd_sc_hd__clkbuf_1
X_4439_ _4519_/A _4547_/B vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__nand2_1
XFILLER_120_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6843__103 vssd1 vssd1 vccd1 vccd1 _6843__103/HI _6952_/A sky130_fd_sc_hd__conb_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6109_ _6760_/Q _6106_/X _6108_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6110_/B sky130_fd_sc_hd__a22o_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3810_ _3810_/A _3810_/B vssd1 vssd1 vccd1 vccd1 _3811_/B sky130_fd_sc_hd__nand2_1
X_4790_ _4790_/A vssd1 vssd1 vccd1 vccd1 _6460_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_29 _3325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3741_ _3741_/A _3741_/B _3741_/C vssd1 vssd1 vccd1 vccd1 _3745_/B sky130_fd_sc_hd__nand3_1
XANTENNA_18 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3672_ _3669_/X _3670_/Y _3671_/X _3629_/A vssd1 vssd1 vccd1 vccd1 _3674_/A sky130_fd_sc_hd__o211a_1
X_6460_ _6789_/CLK _6460_/D vssd1 vssd1 vccd1 vccd1 _6460_/Q sky130_fd_sc_hd__dfxtp_1
X_5411_ _3349_/X _5406_/X _5331_/X vssd1 vssd1 vccd1 vccd1 _6646_/D sky130_fd_sc_hd__o21a_1
X_6391_ _6795_/CLK _6391_/D vssd1 vssd1 vccd1 vccd1 _6391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5342_ _6207_/A vssd1 vssd1 vccd1 vccd1 _5342_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5273_ _5273_/A vssd1 vssd1 vccd1 vccd1 _5282_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4224_ _4224_/A vssd1 vssd1 vccd1 vccd1 _6370_/D sky130_fd_sc_hd__clkbuf_1
X_4155_ _4155_/A _4155_/B vssd1 vssd1 vccd1 vccd1 _4157_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4086_ _4086_/A _4086_/B vssd1 vssd1 vccd1 vccd1 _4087_/B sky130_fd_sc_hd__nor2_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4988_ _4988_/A vssd1 vssd1 vccd1 vccd1 _6545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3939_ _4013_/A _4268_/A vssd1 vssd1 vccd1 vccd1 _3940_/B sky130_fd_sc_hd__nand2_1
X_6727_ _6799_/CLK _6727_/D vssd1 vssd1 vccd1 vccd1 _6727_/Q sky130_fd_sc_hd__dfxtp_1
X_6658_ _6795_/CLK _6658_/D vssd1 vssd1 vccd1 vccd1 _6658_/Q sky130_fd_sc_hd__dfxtp_1
X_5609_ _6680_/Q _5601_/X _5606_/X _5608_/X _5591_/X vssd1 vssd1 vccd1 vccd1 _6680_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6589_ _6667_/CLK _6589_/D vssd1 vssd1 vccd1 vccd1 _6589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput16 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _3330_/A sky130_fd_sc_hd__buf_2
Xinput27 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_4
Xinput38 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_2
Xinput49 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5960_ _6734_/Q _5946_/X _5958_/X _5959_/X vssd1 vssd1 vccd1 vccd1 _6734_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4911_ _4911_/A vssd1 vssd1 vccd1 vccd1 _6525_/D sky130_fd_sc_hd__clkbuf_1
X_5891_ _5920_/A vssd1 vssd1 vccd1 vccd1 _5891_/X sky130_fd_sc_hd__clkbuf_2
X_4842_ _4842_/A vssd1 vssd1 vccd1 vccd1 _6483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4773_ _4773_/A vssd1 vssd1 vccd1 vccd1 _6452_/D sky130_fd_sc_hd__clkbuf_1
X_6512_ _6522_/CLK _6512_/D vssd1 vssd1 vccd1 vccd1 _6512_/Q sky130_fd_sc_hd__dfxtp_1
X_3724_ _3724_/A _3765_/B _3724_/C vssd1 vssd1 vccd1 vccd1 _3769_/A sky130_fd_sc_hd__and3_1
XFILLER_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6443_ _6795_/CLK _6443_/D vssd1 vssd1 vccd1 vccd1 _6443_/Q sky130_fd_sc_hd__dfxtp_1
X_3655_ _3656_/B _3656_/C _3656_/A vssd1 vssd1 vccd1 vccd1 _3679_/B sky130_fd_sc_hd__a21o_1
X_6374_ _6795_/CLK _6374_/D vssd1 vssd1 vccd1 vccd1 _6374_/Q sky130_fd_sc_hd__dfxtp_1
X_3586_ _3586_/A _3586_/B _3586_/C vssd1 vssd1 vccd1 vccd1 _3614_/A sky130_fd_sc_hd__nor3_2
XFILLER_102_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5325_ _5502_/B _5964_/C _3637_/A vssd1 vssd1 vccd1 vccd1 _5325_/Y sky130_fd_sc_hd__a21oi_1
X_5256_ _6594_/Q _5260_/B vssd1 vssd1 vccd1 vccd1 _5257_/A sky130_fd_sc_hd__and2_1
X_4207_ _4186_/B _4207_/B vssd1 vssd1 vccd1 vccd1 _4207_/X sky130_fd_sc_hd__and2b_1
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5187_ _6920_/A _5209_/B vssd1 vssd1 vccd1 vccd1 _5191_/B sky130_fd_sc_hd__or2_1
XFILLER_95_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4138_ _4169_/B _4169_/C _4169_/A vssd1 vssd1 vccd1 vccd1 _4140_/A sky130_fd_sc_hd__a21o_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4069_ _4067_/X _4026_/A _4065_/Y _4066_/X vssd1 vssd1 vccd1 vccd1 _4069_/X sky130_fd_sc_hd__a211o_1
XFILLER_44_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3440_ _5214_/B vssd1 vssd1 vccd1 vccd1 _3879_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3371_ _6495_/Q _3370_/B _6496_/Q vssd1 vssd1 vccd1 vccd1 _3372_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5110_ _5081_/X _5108_/X _5109_/X _5088_/X vssd1 vssd1 vccd1 vccd1 _5110_/X sky130_fd_sc_hd__a31o_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6090_ _6110_/A _6090_/B vssd1 vssd1 vccd1 vccd1 _6091_/A sky130_fd_sc_hd__and2_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A vssd1 vssd1 vccd1 vccd1 _5041_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6992_ _6992_/A _3298_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5943_ _6489_/Q _5957_/B _5943_/C vssd1 vssd1 vccd1 vccd1 _5943_/X sky130_fd_sc_hd__and3_1
X_5874_ _5941_/A vssd1 vssd1 vccd1 vccd1 _5874_/X sky130_fd_sc_hd__buf_2
X_4825_ _4847_/A vssd1 vssd1 vccd1 vccd1 _4834_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_21_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4756_ _6397_/Q _4756_/B vssd1 vssd1 vccd1 vccd1 _4757_/A sky130_fd_sc_hd__and2_1
X_3707_ _3639_/A _5214_/A _3663_/B _3706_/X vssd1 vssd1 vccd1 vccd1 _3709_/A sky130_fd_sc_hd__a31o_1
X_4687_ _4687_/A vssd1 vssd1 vccd1 vccd1 _6414_/D sky130_fd_sc_hd__clkbuf_1
X_6426_ _6763_/CLK _6426_/D vssd1 vssd1 vccd1 vccd1 _6426_/Q sky130_fd_sc_hd__dfxtp_1
X_3638_ _3706_/A _5214_/C _3638_/C vssd1 vssd1 vccd1 vccd1 _3638_/X sky130_fd_sc_hd__and3_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3569_ _3706_/A _5217_/A _3569_/C vssd1 vssd1 vccd1 vccd1 _3569_/X sky130_fd_sc_hd__and3_1
X_6357_ _6763_/CLK _6357_/D vssd1 vssd1 vccd1 vccd1 _6357_/Q sky130_fd_sc_hd__dfxtp_2
X_5308_ _6617_/Q _5346_/B vssd1 vssd1 vccd1 vccd1 _5309_/A sky130_fd_sc_hd__and2_1
X_6288_ _6815_/Q _6230_/X _6287_/Y _6275_/X vssd1 vssd1 vccd1 vccd1 _6815_/D sky130_fd_sc_hd__o211a_1
X_5239_ _5242_/B _5239_/B _5239_/C vssd1 vssd1 vccd1 vccd1 _5240_/A sky130_fd_sc_hd__and3b_1
XFILLER_102_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4610_ _4611_/A _4611_/B vssd1 vssd1 vccd1 vccd1 _4634_/A sky130_fd_sc_hd__or2_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5590_ _6253_/A _5589_/X _5578_/X _5567_/X vssd1 vssd1 vccd1 vccd1 _5590_/X sky130_fd_sc_hd__a31o_1
X_4541_ _4541_/A _4541_/B vssd1 vssd1 vccd1 vccd1 _4541_/Y sky130_fd_sc_hd__nor2_1
X_4472_ _4473_/B _4473_/C _4473_/A vssd1 vssd1 vccd1 vccd1 _4475_/A sky130_fd_sc_hd__a21o_1
X_6211_ _6270_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6211_/X sky130_fd_sc_hd__or2_1
X_3423_ _3423_/A vssd1 vssd1 vccd1 vccd1 _6299_/D sky130_fd_sc_hd__clkbuf_1
X_6142_ _6169_/A vssd1 vssd1 vccd1 vccd1 _6142_/X sky130_fd_sc_hd__clkbuf_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3354_ _6224_/B vssd1 vssd1 vccd1 vccd1 _6102_/A sky130_fd_sc_hd__buf_2
XFILLER_58_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3286_/A vssd1 vssd1 vccd1 vccd1 _3285_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6073_ _6084_/A _6073_/B vssd1 vssd1 vccd1 vccd1 _6074_/A sky130_fd_sc_hd__and2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _6537_/Q _6535_/Q vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__nor2_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6975_ _6975_/A _3278_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
X_5926_ _5602_/X _5919_/X _5920_/X _5912_/X _6728_/Q vssd1 vssd1 vccd1 vccd1 _5926_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_41_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5857_ _6491_/Q _5840_/X _5856_/X _5836_/X _5843_/X vssd1 vssd1 vccd1 vccd1 _5857_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4808_ _6420_/Q _4812_/B vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__and2_1
X_5788_ _5843_/A vssd1 vssd1 vccd1 vccd1 _5788_/X sky130_fd_sc_hd__clkbuf_2
X_4739_ _4739_/A vssd1 vssd1 vccd1 vccd1 _6437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6409_ _6789_/CLK _6409_/D vssd1 vssd1 vccd1 vccd1 _6409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6760_ _6763_/CLK _6760_/D vssd1 vssd1 vccd1 vccd1 _6760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5711_ _6240_/A _5678_/X _5680_/X _5710_/X _5695_/X vssd1 vssd1 vccd1 vccd1 _5711_/X
+ sky130_fd_sc_hd__a221o_1
X_3972_ _4121_/A _4121_/B _4076_/C _6352_/Q vssd1 vssd1 vccd1 vccd1 _3972_/X sky130_fd_sc_hd__and4_1
X_6691_ _6789_/CLK _6691_/D vssd1 vssd1 vccd1 vccd1 _6691_/Q sky130_fd_sc_hd__dfxtp_1
X_5642_ _6474_/Q vssd1 vssd1 vccd1 vccd1 _5642_/X sky130_fd_sc_hd__buf_2
X_5573_ _5669_/S vssd1 vssd1 vccd1 vccd1 _5612_/S sky130_fd_sc_hd__clkbuf_2
X_4524_ _4524_/A _4524_/B _4524_/C vssd1 vssd1 vccd1 vccd1 _4540_/B sky130_fd_sc_hd__nand3_2
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4455_ _4455_/A _4455_/B _4455_/C vssd1 vssd1 vccd1 vccd1 _4455_/X sky130_fd_sc_hd__and3_2
X_3406_ _3486_/A vssd1 vssd1 vccd1 vccd1 _3499_/S sky130_fd_sc_hd__buf_4
X_4386_ _4382_/X _4383_/X _4385_/X vssd1 vssd1 vccd1 vccd1 _6387_/D sky130_fd_sc_hd__a21oi_1
XFILLER_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3337_ _3377_/A vssd1 vssd1 vccd1 vccd1 _5284_/A sky130_fd_sc_hd__buf_2
XFILLER_86_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6125_ _6125_/A vssd1 vssd1 vccd1 vccd1 _6763_/D sky130_fd_sc_hd__clkbuf_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6056_ _6493_/Q _6056_/B _6056_/C vssd1 vssd1 vccd1 vccd1 _6056_/X sky130_fd_sc_hd__and3_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _3268_/A vssd1 vssd1 vccd1 vccd1 _3268_/Y sky130_fd_sc_hd__inv_2
X_5007_ _5006_/Y hold2/A _6330_/D vssd1 vssd1 vccd1 vccd1 _6552_/D sky130_fd_sc_hd__a21o_1
X_3199_ _3200_/A vssd1 vssd1 vccd1 vccd1 _3199_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6958_ _6958_/A _3259_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5909_ _6483_/Q _5931_/B _5914_/C vssd1 vssd1 vccd1 vccd1 _5909_/X sky130_fd_sc_hd__and3_1
XFILLER_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4240_ _4235_/A _4239_/Y _4235_/B vssd1 vssd1 vccd1 vccd1 _4240_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4171_ _4220_/A _4220_/C _4170_/Y vssd1 vssd1 vccd1 vccd1 _4172_/B sky130_fd_sc_hd__o21a_1
XFILLER_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6812_ _6532_/Q _6812_/D vssd1 vssd1 vccd1 vccd1 _6812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6743_ _6532_/Q _6743_/D vssd1 vssd1 vccd1 vccd1 _6743_/Q sky130_fd_sc_hd__dfxtp_1
X_3955_ _6067_/A _3955_/B _3988_/B vssd1 vssd1 vccd1 vccd1 _6362_/D sky130_fd_sc_hd__nor3_1
XFILLER_51_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6674_ _6809_/CLK _6674_/D vssd1 vssd1 vccd1 vccd1 _6674_/Q sky130_fd_sc_hd__dfxtp_1
X_5625_ _5619_/X _5582_/X _5620_/X _5624_/X vssd1 vssd1 vccd1 vccd1 _5625_/X sky130_fd_sc_hd__o211a_1
X_3886_ _6350_/Q vssd1 vssd1 vccd1 vccd1 _4039_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5556_ _5552_/X _5525_/X _5505_/X _5555_/X vssd1 vssd1 vccd1 vccd1 _5556_/X sky130_fd_sc_hd__o211a_1
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4507_ _4505_/X _4615_/A _3637_/A vssd1 vssd1 vccd1 vccd1 _4507_/Y sky130_fd_sc_hd__a21oi_1
X_5487_ _5490_/A _5487_/B vssd1 vssd1 vccd1 vccd1 _5488_/A sky130_fd_sc_hd__and2_1
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4438_ _4437_/B _4437_/C _4437_/A vssd1 vssd1 vccd1 vccd1 _4445_/C sky130_fd_sc_hd__a21o_1
X_6882__142 vssd1 vssd1 vccd1 vccd1 _6882__142/HI _6991_/A sky130_fd_sc_hd__conb_1
X_4369_ _4519_/A _4371_/B _4366_/Y _4368_/X vssd1 vssd1 vccd1 vccd1 _4369_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6108_ _6470_/Q _6107_/X _6096_/X _6087_/X _6486_/Q vssd1 vssd1 vccd1 vccd1 _6108_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6039_ _6748_/Q _5642_/X _6044_/S vssd1 vssd1 vccd1 vccd1 _6039_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_19 _5008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3740_ _3737_/Y _3738_/X _3703_/B _3703_/Y vssd1 vssd1 vccd1 vccd1 _3741_/C sky130_fd_sc_hd__o211ai_2
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3671_ _3671_/A _3671_/B _3671_/C vssd1 vssd1 vccd1 vccd1 _3671_/X sky130_fd_sc_hd__or3_1
X_5410_ _5410_/A vssd1 vssd1 vccd1 vccd1 _6645_/D sky130_fd_sc_hd__clkbuf_1
X_6390_ _6795_/CLK _6390_/D vssd1 vssd1 vccd1 vccd1 _6390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5341_ _5870_/A _6143_/A vssd1 vssd1 vccd1 vccd1 _6207_/A sky130_fd_sc_hd__nor2_2
X_6866__126 vssd1 vssd1 vccd1 vccd1 _6866__126/HI _6975_/A sky130_fd_sc_hd__conb_1
X_5272_ _5272_/A vssd1 vssd1 vccd1 vccd1 _6601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4223_ _4221_/X _4223_/B vssd1 vssd1 vccd1 vccd1 _4224_/A sky130_fd_sc_hd__and2b_1
X_4154_ _4154_/A _4154_/B vssd1 vssd1 vccd1 vccd1 _4155_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4085_ _4147_/A _4085_/B _6354_/Q _4180_/D vssd1 vssd1 vccd1 vccd1 _4086_/B sky130_fd_sc_hd__and4_1
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4987_ _5129_/A _4987_/B _4987_/C vssd1 vssd1 vccd1 vccd1 _4988_/A sky130_fd_sc_hd__and3_1
X_6726_ _6809_/CLK _6726_/D vssd1 vssd1 vccd1 vccd1 _6726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3938_ _4116_/B vssd1 vssd1 vccd1 vccd1 _4268_/A sky130_fd_sc_hd__buf_2
X_6657_ _6795_/CLK _6657_/D vssd1 vssd1 vccd1 vccd1 _6657_/Q sky130_fd_sc_hd__dfxtp_1
X_3869_ _5217_/B _6275_/A vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__and2_1
X_6588_ _6667_/CLK _6588_/D vssd1 vssd1 vccd1 vccd1 _6588_/Q sky130_fd_sc_hd__dfxtp_1
X_5608_ _6260_/A _5589_/X _5578_/X _5567_/X vssd1 vssd1 vccd1 vccd1 _5608_/X sky130_fd_sc_hd__a31o_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5539_ _6233_/A _5534_/X _6286_/B _5538_/X vssd1 vssd1 vccd1 vccd1 _5539_/X sky130_fd_sc_hd__a31o_1
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _3326_/C sky130_fd_sc_hd__clkbuf_4
Xinput17 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 _3330_/D sky130_fd_sc_hd__buf_2
Xinput39 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_2
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4910_ _4909_/X _6525_/Q _4910_/S vssd1 vssd1 vccd1 vccd1 _4911_/A sky130_fd_sc_hd__mux2_1
X_5890_ _5890_/A vssd1 vssd1 vccd1 vccd1 _5920_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4841_ _6435_/Q _4845_/B vssd1 vssd1 vccd1 vccd1 _4842_/A sky130_fd_sc_hd__and2_1
X_4772_ _6404_/Q _4778_/B vssd1 vssd1 vccd1 vccd1 _4773_/A sky130_fd_sc_hd__and2_1
X_6511_ _6522_/CLK _6511_/D vssd1 vssd1 vccd1 vccd1 _6511_/Q sky130_fd_sc_hd__dfxtp_1
X_3723_ _3684_/A _3684_/B _3684_/C vssd1 vssd1 vccd1 vccd1 _3724_/C sky130_fd_sc_hd__a21bo_1
XFILLER_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6442_ _6795_/CLK _6442_/D vssd1 vssd1 vccd1 vccd1 _6442_/Q sky130_fd_sc_hd__dfxtp_1
X_3654_ _3698_/A _3698_/B vssd1 vssd1 vccd1 vccd1 _3656_/A sky130_fd_sc_hd__xor2_1
X_6373_ _6795_/CLK _6373_/D vssd1 vssd1 vccd1 vccd1 _6373_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_3585_ _3585_/A _3585_/B _3585_/C vssd1 vssd1 vccd1 vccd1 _3586_/C sky130_fd_sc_hd__and3_1
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5324_ _5337_/B vssd1 vssd1 vccd1 vccd1 _5964_/C sky130_fd_sc_hd__clkbuf_2
X_5255_ _5255_/A vssd1 vssd1 vccd1 vccd1 _6593_/D sky130_fd_sc_hd__clkbuf_1
X_4206_ _4243_/A _4206_/B vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__or2_1
X_5186_ _5186_/A vssd1 vssd1 vccd1 vccd1 _5209_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _4106_/A _4106_/C _4106_/B vssd1 vssd1 vccd1 vccd1 _4169_/A sky130_fd_sc_hd__a21bo_1
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4068_ _4065_/Y _4066_/X _4067_/X _4026_/A vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__o211a_1
XFILLER_83_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6709_ _6809_/CLK _6709_/D vssd1 vssd1 vccd1 vccd1 _6709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3370_ _6495_/Q _3370_/B vssd1 vssd1 vccd1 vccd1 _6495_/D sky130_fd_sc_hd__xor2_1
XFILLER_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5040_ _6896_/A _4945_/X _5039_/X _5034_/X vssd1 vssd1 vccd1 vccd1 _6558_/D sky130_fd_sc_hd__o211a_1
XFILLER_78_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6991_ _6991_/A _3297_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
XFILLER_65_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5942_ _5630_/X _5919_/X _5920_/X _5961_/B _6731_/Q vssd1 vssd1 vccd1 vccd1 _5942_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5873_ _5873_/A _5890_/A vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4824_ _4824_/A vssd1 vssd1 vccd1 vccd1 _6475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4755_ _4755_/A vssd1 vssd1 vccd1 vccd1 _6444_/D sky130_fd_sc_hd__clkbuf_1
X_3706_ _3706_/A _5214_/B _3706_/C vssd1 vssd1 vccd1 vccd1 _3706_/X sky130_fd_sc_hd__and3_1
XFILLER_107_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4686_ _6358_/Q _4688_/B vssd1 vssd1 vccd1 vccd1 _4687_/A sky130_fd_sc_hd__and2_1
X_3637_ _3637_/A vssd1 vssd1 vccd1 vccd1 _4990_/A sky130_fd_sc_hd__buf_4
X_6425_ _6763_/CLK _6425_/D vssd1 vssd1 vccd1 vccd1 _6425_/Q sky130_fd_sc_hd__dfxtp_1
X_6356_ _6763_/CLK _6356_/D vssd1 vssd1 vccd1 vccd1 _6356_/Q sky130_fd_sc_hd__dfxtp_1
X_3568_ _3568_/A vssd1 vssd1 vccd1 vccd1 _3593_/A sky130_fd_sc_hd__inv_2
XFILLER_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5307_ _5374_/A vssd1 vssd1 vccd1 vccd1 _5346_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3499_ _6327_/Q _6531_/Q _3499_/S vssd1 vssd1 vccd1 vccd1 _3500_/A sky130_fd_sc_hd__mux2_1
X_6287_ _6248_/A _6286_/Y _6267_/A vssd1 vssd1 vccd1 vccd1 _6287_/Y sky130_fd_sc_hd__o21ai_1
X_5238_ _6587_/Q _5238_/B vssd1 vssd1 vccd1 vccd1 _5239_/C sky130_fd_sc_hd__or2_1
XFILLER_84_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5169_ _5169_/A vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4540_ _4540_/A _4540_/B _4540_/C vssd1 vssd1 vccd1 vccd1 _4540_/Y sky130_fd_sc_hd__nand3_1
X_4471_ _6669_/Q _6377_/Q vssd1 vssd1 vccd1 vccd1 _4473_/A sky130_fd_sc_hd__and2_1
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6210_ _6793_/Q _6207_/X _6209_/X _6203_/X vssd1 vssd1 vccd1 vccd1 _6793_/D sky130_fd_sc_hd__o211a_1
X_3422_ _5217_/A _6503_/Q _3427_/S vssd1 vssd1 vccd1 vccd1 _3423_/A sky130_fd_sc_hd__mux2_1
X_6141_ _6143_/A _6143_/B vssd1 vssd1 vccd1 vccd1 _6169_/A sky130_fd_sc_hd__nor2_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3353_ _3349_/X _5406_/A _5406_/B _3352_/X vssd1 vssd1 vccd1 vccd1 _6224_/B sky130_fd_sc_hd__a31oi_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6072_ _6753_/Q _6061_/X _6071_/X _5824_/A vssd1 vssd1 vccd1 vccd1 _6073_/B sky130_fd_sc_hd__a22o_1
X_3284_ _3286_/A vssd1 vssd1 vccd1 vccd1 _3284_/Y sky130_fd_sc_hd__inv_2
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5023_ _5043_/A _5023_/B vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__or2_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6974_ _6974_/A _3277_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
XFILLER_110_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _6727_/Q _5918_/X _5924_/X _5904_/X vssd1 vssd1 vccd1 vccd1 _6727_/D sky130_fd_sc_hd__o211a_1
X_5856_ _5651_/X _5855_/X _5860_/S vssd1 vssd1 vccd1 vccd1 _5856_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4807_ _4807_/A vssd1 vssd1 vccd1 vccd1 _6467_/D sky130_fd_sc_hd__clkbuf_1
X_5787_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5787_/X sky130_fd_sc_hd__clkbuf_2
X_4738_ _6389_/Q _4744_/B vssd1 vssd1 vccd1 vccd1 _4739_/A sky130_fd_sc_hd__and2_1
XFILLER_107_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4669_ _6342_/Q _4677_/B vssd1 vssd1 vccd1 vccd1 _4670_/A sky130_fd_sc_hd__and2_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6408_ _6789_/CLK _6408_/D vssd1 vssd1 vccd1 vccd1 _6408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6339_ _6789_/CLK _6339_/D vssd1 vssd1 vccd1 vccd1 _6339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3971_ _6660_/Q vssd1 vssd1 vccd1 vccd1 _4121_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5710_ _5552_/X _5709_/X _5721_/S vssd1 vssd1 vccd1 vccd1 _5710_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6690_ _6809_/CLK _6690_/D vssd1 vssd1 vccd1 vccd1 _6690_/Q sky130_fd_sc_hd__dfxtp_1
X_5641_ _6683_/Q _5601_/X _5636_/X _5639_/X _5640_/X vssd1 vssd1 vccd1 vccd1 _6683_/D
+ sky130_fd_sc_hd__o221a_1
X_5572_ _6451_/Q _5603_/B vssd1 vssd1 vccd1 vccd1 _5572_/X sky130_fd_sc_hd__and2_2
X_4523_ _4483_/A _4483_/C _4483_/B vssd1 vssd1 vccd1 vccd1 _4524_/C sky130_fd_sc_hd__a21bo_1
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4454_ _4455_/B _4455_/C _4455_/A vssd1 vssd1 vccd1 vccd1 _4454_/Y sky130_fd_sc_hd__a21oi_2
X_3405_ _3405_/A _6495_/Q _3370_/B vssd1 vssd1 vccd1 vccd1 _3486_/A sky130_fd_sc_hd__nor3b_2
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4385_ _4385_/A _4385_/B vssd1 vssd1 vccd1 vccd1 _4385_/X sky130_fd_sc_hd__or2_1
X_3336_ _4980_/B _4993_/A _5017_/A _6333_/Q vssd1 vssd1 vccd1 vccd1 _3336_/X sky130_fd_sc_hd__and4b_1
X_6124_ _6132_/A _6124_/B vssd1 vssd1 vccd1 vccd1 _6125_/A sky130_fd_sc_hd__and2_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6055_ _5519_/X _6053_/X _6054_/X vssd1 vssd1 vccd1 vccd1 _6055_/X sky130_fd_sc_hd__o21a_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3268_/A vssd1 vssd1 vccd1 vccd1 _3267_/Y sky130_fd_sc_hd__inv_2
X_5006_ _6330_/Q vssd1 vssd1 vccd1 vccd1 _5006_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3198_ _3200_/A vssd1 vssd1 vccd1 vccd1 _3198_/Y sky130_fd_sc_hd__inv_2
X_6957_ _6957_/A _3258_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5908_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5931_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5839_ _6713_/Q _5825_/X _5837_/X _5838_/X vssd1 vssd1 vccd1 vccd1 _6713_/D sky130_fd_sc_hd__o211a_1
XFILLER_6_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4170_ _4168_/A _4169_/X _4140_/A vssd1 vssd1 vccd1 vccd1 _4170_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6811_ _6532_/Q _6811_/D vssd1 vssd1 vccd1 vccd1 _6811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6742_ _6799_/CLK _6742_/D vssd1 vssd1 vccd1 vccd1 _6742_/Q sky130_fd_sc_hd__dfxtp_1
X_3954_ _3953_/A _3953_/B _3953_/C vssd1 vssd1 vccd1 vccd1 _3988_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6673_ _6809_/CLK _6673_/D vssd1 vssd1 vccd1 vccd1 _6673_/Q sky130_fd_sc_hd__dfxtp_1
X_3885_ _4056_/A vssd1 vssd1 vccd1 vccd1 _3889_/A sky130_fd_sc_hd__clkbuf_2
X_5624_ _5624_/A _5624_/B vssd1 vssd1 vccd1 vccd1 _5624_/X sky130_fd_sc_hd__or2_1
X_5555_ _5575_/A _5555_/B vssd1 vssd1 vccd1 vccd1 _5555_/X sky130_fd_sc_hd__or2_1
X_4506_ _4463_/A _4463_/B _4462_/B _4460_/X vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__a31o_1
X_5486_ _6316_/Q _4574_/A _5496_/S vssd1 vssd1 vccd1 vccd1 _5487_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4437_ _4437_/A _4437_/B _4437_/C vssd1 vssd1 vccd1 vccd1 _4445_/B sky130_fd_sc_hd__nand3_1
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4368_ _4368_/A _4368_/B _4433_/D _4510_/C vssd1 vssd1 vccd1 vccd1 _4368_/X sky130_fd_sc_hd__and4_1
X_6107_ _6107_/A vssd1 vssd1 vccd1 vccd1 _6107_/X sky130_fd_sc_hd__clkbuf_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3377_/A vssd1 vssd1 vccd1 vccd1 _3632_/A sky130_fd_sc_hd__clkinv_2
X_4299_ _4451_/A _4296_/C _4333_/B _4407_/A vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__a22o_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6038_ _6747_/Q _6011_/X _6037_/X _6027_/X vssd1 vssd1 vccd1 vccd1 _6747_/D sky130_fd_sc_hd__o211a_1
XFILLER_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6504_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_82_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3670_ _3667_/X _3668_/Y _3638_/X _3639_/X vssd1 vssd1 vccd1 vccd1 _3670_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5340_ _5335_/X _6192_/B _6330_/D vssd1 vssd1 vccd1 vccd1 _6622_/D sky130_fd_sc_hd__a21o_1
X_5271_ _6601_/Q _5271_/B vssd1 vssd1 vccd1 vccd1 _5272_/A sky130_fd_sc_hd__and2_1
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4222_ _4219_/X _4220_/X _4217_/Y vssd1 vssd1 vccd1 vccd1 _4223_/B sky130_fd_sc_hd__a21o_1
X_4153_ _4153_/A _4153_/B _4153_/C _6354_/Q vssd1 vssd1 vccd1 vccd1 _4154_/B sky130_fd_sc_hd__and4_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4084_ _4147_/A _4180_/C _4180_/D _4085_/B vssd1 vssd1 vccd1 vccd1 _4086_/A sky130_fd_sc_hd__a22oi_1
XFILLER_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4986_ _6545_/Q _4986_/B vssd1 vssd1 vccd1 vccd1 _4987_/C sky130_fd_sc_hd__nand2_1
XFILLER_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3937_ _6354_/Q vssd1 vssd1 vccd1 vccd1 _4116_/B sky130_fd_sc_hd__clkbuf_2
X_6725_ _6809_/CLK _6725_/D vssd1 vssd1 vccd1 vccd1 _6725_/Q sky130_fd_sc_hd__dfxtp_1
X_6656_ _6795_/CLK _6656_/D vssd1 vssd1 vccd1 vccd1 _6656_/Q sky130_fd_sc_hd__dfxtp_1
X_3868_ _3868_/A vssd1 vssd1 vccd1 vccd1 _6351_/D sky130_fd_sc_hd__clkbuf_1
X_6587_ _6667_/CLK _6587_/D vssd1 vssd1 vccd1 vccd1 _6587_/Q sky130_fd_sc_hd__dfxtp_1
X_5607_ _6486_/Q vssd1 vssd1 vccd1 vccd1 _6260_/A sky130_fd_sc_hd__clkbuf_4
X_3799_ _3797_/Y _3767_/B _3798_/X vssd1 vssd1 vccd1 vccd1 _3820_/B sky130_fd_sc_hd__a21bo_1
X_5538_ _5843_/A vssd1 vssd1 vccd1 vccd1 _5538_/X sky130_fd_sc_hd__buf_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5469_ _5469_/A vssd1 vssd1 vccd1 vccd1 _5483_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_87_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _3330_/C sky130_fd_sc_hd__buf_4
Xinput29 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _3325_/B sky130_fd_sc_hd__buf_4
X_6889__149 vssd1 vssd1 vccd1 vccd1 _6889__149/HI _6998_/A sky130_fd_sc_hd__conb_1
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4840_ _4840_/A vssd1 vssd1 vccd1 vccd1 _6482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6510_ _6523_/CLK _6510_/D vssd1 vssd1 vccd1 vccd1 _6510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4771_ _4771_/A vssd1 vssd1 vccd1 vccd1 _6451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3722_ _3757_/A _3722_/B _3722_/C _3765_/A vssd1 vssd1 vccd1 vccd1 _3765_/B sky130_fd_sc_hd__nand4_1
X_6441_ _6795_/CLK _6441_/D vssd1 vssd1 vccd1 vccd1 _6441_/Q sky130_fd_sc_hd__dfxtp_1
X_3653_ _3653_/A _3653_/B vssd1 vssd1 vccd1 vccd1 _3698_/B sky130_fd_sc_hd__or2_1
X_6372_ _6795_/CLK _6372_/D vssd1 vssd1 vccd1 vccd1 _6372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5323_ _5518_/A _5499_/B vssd1 vssd1 vccd1 vccd1 _5337_/B sky130_fd_sc_hd__nor2_1
X_3584_ _3585_/B _3585_/C _3585_/A vssd1 vssd1 vccd1 vccd1 _3586_/B sky130_fd_sc_hd__a21oi_1
X_5254_ _6593_/Q _5260_/B vssd1 vssd1 vccd1 vccd1 _5255_/A sky130_fd_sc_hd__and2_1
X_5185_ _5185_/A vssd1 vssd1 vccd1 vccd1 _6581_/D sky130_fd_sc_hd__clkbuf_1
X_4205_ _4205_/A _4205_/B _4205_/C vssd1 vssd1 vccd1 vccd1 _4206_/B sky130_fd_sc_hd__nor3_1
XFILLER_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4136_ _4135_/B _4135_/C _4135_/A vssd1 vssd1 vccd1 vccd1 _4169_/C sky130_fd_sc_hd__a21o_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4067_ _4067_/A _4067_/B _4067_/C vssd1 vssd1 vccd1 vccd1 _4067_/X sky130_fd_sc_hd__or3_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4969_ _6540_/Q _6539_/Q _4969_/C vssd1 vssd1 vccd1 vccd1 _4972_/B sky130_fd_sc_hd__and3_1
X_6708_ _6809_/CLK _6708_/D vssd1 vssd1 vccd1 vccd1 _6708_/Q sky130_fd_sc_hd__dfxtp_1
X_6639_ _6532_/Q _6639_/D vssd1 vssd1 vccd1 vccd1 _6639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6990_ _6990_/A _3296_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
XFILLER_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5941_ _5941_/A vssd1 vssd1 vccd1 vccd1 _5961_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5872_ _5872_/A _5872_/B vssd1 vssd1 vccd1 vccd1 _5890_/A sky130_fd_sc_hd__nor2_2
XFILLER_80_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4823_ _6427_/Q _4823_/B vssd1 vssd1 vccd1 vccd1 _4824_/A sky130_fd_sc_hd__and2_1
XFILLER_21_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4754_ _6396_/Q _4756_/B vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__and2_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ _3702_/X _3703_/Y _3679_/X _3665_/X vssd1 vssd1 vccd1 vccd1 _3709_/C sky130_fd_sc_hd__a211o_1
X_4685_ _4685_/A vssd1 vssd1 vccd1 vccd1 _6413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3636_ _3636_/A vssd1 vssd1 vccd1 vccd1 _3637_/A sky130_fd_sc_hd__clkbuf_4
X_6424_ _6763_/CLK _6424_/D vssd1 vssd1 vccd1 vccd1 _6424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6355_ _6763_/CLK _6355_/D vssd1 vssd1 vccd1 vccd1 _6355_/Q sky130_fd_sc_hd__dfxtp_1
X_3567_ _6067_/A _3567_/B _3593_/B vssd1 vssd1 vccd1 vccd1 _6338_/D sky130_fd_sc_hd__nor3_1
XFILLER_115_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5306_ _5306_/A vssd1 vssd1 vccd1 vccd1 _6616_/D sky130_fd_sc_hd__clkbuf_1
X_6286_ _6286_/A _6286_/B vssd1 vssd1 vccd1 vccd1 _6286_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5237_ _6587_/Q _5238_/B vssd1 vssd1 vccd1 vccd1 _5242_/B sky130_fd_sc_hd__and2_1
XFILLER_102_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3498_ _3498_/A vssd1 vssd1 vccd1 vccd1 _6326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5168_ _6917_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5172_/B sky130_fd_sc_hd__or2_1
XFILLER_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5099_ _5081_/X _5097_/X _5098_/X _5088_/X vssd1 vssd1 vccd1 vccd1 _5099_/X sky130_fd_sc_hd__a31o_1
XFILLER_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4119_ _4118_/A _4156_/B _4118_/C vssd1 vssd1 vccd1 vccd1 _4146_/B sky130_fd_sc_hd__a21oi_1
XFILLER_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4470_ _6671_/Q _4510_/B _6375_/Q _4510_/C vssd1 vssd1 vccd1 vccd1 _4473_/C sky130_fd_sc_hd__nand4_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3421_ _3762_/D vssd1 vssd1 vccd1 vccd1 _5217_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3352_ _6647_/Q _6329_/Q vssd1 vssd1 vccd1 vccd1 _3352_/X sky130_fd_sc_hd__or2b_1
X_6140_ _6061_/X _6138_/X _6139_/X _6051_/X vssd1 vssd1 vccd1 vccd1 _6767_/D sky130_fd_sc_hd__o211a_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _5524_/X _5947_/X _6070_/X _6138_/S _6479_/Q vssd1 vssd1 vccd1 vccd1 _6071_/X
+ sky130_fd_sc_hd__a32o_1
X_3283_ _3286_/A vssd1 vssd1 vccd1 vccd1 _3283_/Y sky130_fd_sc_hd__inv_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5022_ _6673_/Q _6705_/Q _6737_/Q _6769_/Q _5012_/X _5014_/X vssd1 vssd1 vccd1 vccd1
+ _5023_/B sky130_fd_sc_hd__mux4_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6973_ _6973_/A _3276_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
XFILLER_80_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5924_ _5906_/X _5921_/X _5923_/X _5915_/X vssd1 vssd1 vccd1 vccd1 _5924_/X sky130_fd_sc_hd__a211o_1
X_5855_ _6717_/Q _5652_/X _5859_/S vssd1 vssd1 vccd1 vccd1 _5855_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4806_ _6419_/Q _4812_/B vssd1 vssd1 vccd1 vccd1 _4807_/A sky130_fd_sc_hd__and2_1
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6584_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_5786_ _6268_/A _5876_/B _5786_/C _6224_/C vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__and4b_2
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4737_ _4737_/A vssd1 vssd1 vccd1 vccd1 _6436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4668_ _4679_/A vssd1 vssd1 vccd1 vccd1 _4677_/B sky130_fd_sc_hd__clkbuf_1
X_6407_ _6789_/CLK _6407_/D vssd1 vssd1 vccd1 vccd1 _6407_/Q sky130_fd_sc_hd__dfxtp_1
X_3619_ _3638_/C _3619_/B vssd1 vssd1 vccd1 vccd1 _3639_/C sky130_fd_sc_hd__xnor2_1
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4599_ _4600_/A _4600_/B _4600_/C vssd1 vssd1 vccd1 vccd1 _4638_/A sky130_fd_sc_hd__o21a_1
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6338_ _6789_/CLK _6338_/D vssd1 vssd1 vccd1 vccd1 _6338_/Q sky130_fd_sc_hd__dfxtp_1
X_6269_ _6269_/A vssd1 vssd1 vccd1 vccd1 _6283_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3970_ _3944_/A _4005_/D _3998_/C _4085_/B vssd1 vssd1 vccd1 vccd1 _3970_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5640_ _5707_/A vssd1 vssd1 vccd1 vccd1 _5640_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5571_ _5620_/A vssd1 vssd1 vccd1 vccd1 _5571_/X sky130_fd_sc_hd__clkbuf_2
X_4522_ _4557_/A _4542_/B _4520_/X vssd1 vssd1 vccd1 vccd1 _4524_/B sky130_fd_sc_hd__or3b_1
X_4453_ _4453_/A _4453_/B vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__xnor2_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3404_ _5217_/D vssd1 vssd1 vccd1 vccd1 _3865_/A sky130_fd_sc_hd__clkbuf_2
X_4384_ _4349_/A _4350_/A _4348_/A _4348_/B _4381_/B vssd1 vssd1 vccd1 vccd1 _4385_/B
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_86_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3335_ _3329_/X _4979_/B _4979_/C _4979_/D vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__and4b_2
X_6123_ _6763_/Q _6106_/X _6122_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6124_/B sky130_fd_sc_hd__a22o_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3268_/A vssd1 vssd1 vccd1 vccd1 _3266_/Y sky130_fd_sc_hd__inv_2
X_6054_ _5667_/X _5990_/S _6751_/Q vssd1 vssd1 vccd1 vccd1 _6054_/X sky130_fd_sc_hd__a21o_1
XFILLER_58_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5005_/A vssd1 vssd1 vccd1 vccd1 _6551_/D sky130_fd_sc_hd__clkbuf_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3197_ _3200_/A vssd1 vssd1 vccd1 vccd1 _3197_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6956_ _6956_/A _3255_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5907_ _5570_/X _5889_/X _5891_/X _5874_/X _6725_/Q vssd1 vssd1 vccd1 vccd1 _5907_/X
+ sky130_fd_sc_hd__a32o_1
X_5838_ _5838_/A vssd1 vssd1 vccd1 vccd1 _5838_/X sky130_fd_sc_hd__clkbuf_2
X_5769_ _6702_/Q _5380_/X _5766_/X _5768_/X _5707_/X vssd1 vssd1 vccd1 vccd1 _6702_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_108_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6810_ _6532_/Q _6810_/D vssd1 vssd1 vccd1 vccd1 _6810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6741_ _6799_/CLK _6741_/D vssd1 vssd1 vccd1 vccd1 _6741_/Q sky130_fd_sc_hd__dfxtp_1
X_3953_ _3953_/A _3953_/B _3953_/C vssd1 vssd1 vccd1 vccd1 _3955_/B sky130_fd_sc_hd__and3_1
XFILLER_51_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6672_ _6809_/CLK _6672_/D vssd1 vssd1 vccd1 vccd1 _6672_/Q sky130_fd_sc_hd__dfxtp_1
X_3884_ _4013_/A vssd1 vssd1 vccd1 vccd1 _4056_/A sky130_fd_sc_hd__clkbuf_2
X_5623_ _6682_/Q _5621_/X _5661_/S vssd1 vssd1 vccd1 vccd1 _5624_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5554_ _6675_/Q _5553_/X _5562_/S vssd1 vssd1 vccd1 vccd1 _5555_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5485_ _5485_/A vssd1 vssd1 vccd1 vccd1 _6667_/D sky130_fd_sc_hd__clkbuf_1
X_4505_ _4566_/A _4566_/B vssd1 vssd1 vccd1 vccd1 _4505_/X sky130_fd_sc_hd__or2_1
X_4436_ _4436_/A _4436_/B _4436_/C vssd1 vssd1 vccd1 vccd1 _4437_/C sky130_fd_sc_hd__nand3_1
XFILLER_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4367_ _6376_/Q vssd1 vssd1 vccd1 vccd1 _4510_/C sky130_fd_sc_hd__clkbuf_2
X_3318_ _3318_/A input2/X vssd1 vssd1 vccd1 vccd1 _3377_/A sky130_fd_sc_hd__nor2_2
XFILLER_59_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6106_ _6106_/A vssd1 vssd1 vccd1 vccd1 _6106_/X sky130_fd_sc_hd__clkbuf_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4298_ _4477_/A vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__clkbuf_2
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3249_ _3249_/A vssd1 vssd1 vccd1 vccd1 _3249_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6037_ _6029_/X _6035_/X _6036_/X vssd1 vssd1 vccd1 vccd1 _6037_/X sky130_fd_sc_hd__a21o_1
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6939_ _6939_/A _3235_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5270_ _5270_/A vssd1 vssd1 vccd1 vccd1 _6600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4221_ _4217_/Y _4219_/X _4220_/X _3636_/A vssd1 vssd1 vccd1 vccd1 _4221_/X sky130_fd_sc_hd__a31o_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4152_ _4153_/A _3998_/D _4180_/C _4180_/B vssd1 vssd1 vccd1 vccd1 _4154_/A sky130_fd_sc_hd__a22oi_2
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4083_ _4083_/A _4183_/B vssd1 vssd1 vccd1 vccd1 _4087_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4985_ _6545_/Q _4986_/B vssd1 vssd1 vccd1 vccd1 _4987_/B sky130_fd_sc_hd__or2_1
X_3936_ _3957_/C _3936_/B vssd1 vssd1 vccd1 vccd1 _3940_/A sky130_fd_sc_hd__xnor2_1
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6724_ _6809_/CLK _6724_/D vssd1 vssd1 vccd1 vccd1 _6724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6655_ _6763_/CLK _6655_/D vssd1 vssd1 vccd1 vccd1 _6655_/Q sky130_fd_sc_hd__dfxtp_2
X_3867_ _5217_/C _6275_/A vssd1 vssd1 vccd1 vccd1 _3868_/A sky130_fd_sc_hd__and2_1
X_6586_ _6586_/CLK _6586_/D vssd1 vssd1 vccd1 vccd1 _6924_/A sky130_fd_sc_hd__dfxtp_1
X_3798_ _3798_/A _3766_/A vssd1 vssd1 vccd1 vccd1 _3798_/X sky130_fd_sc_hd__or2b_1
X_5606_ _5602_/X _5582_/X _5571_/X _5605_/X vssd1 vssd1 vccd1 vccd1 _5606_/X sky130_fd_sc_hd__o211a_1
X_5537_ _6031_/A vssd1 vssd1 vccd1 vccd1 _5843_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5468_ _5468_/A vssd1 vssd1 vccd1 vccd1 _6662_/D sky130_fd_sc_hd__clkbuf_1
X_5399_ _5399_/A vssd1 vssd1 vccd1 vccd1 _6641_/D sky130_fd_sc_hd__clkbuf_1
X_4419_ _4379_/A _4379_/B _4418_/Y vssd1 vssd1 vccd1 vccd1 _4420_/C sky130_fd_sc_hd__a21o_1
XFILLER_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _3333_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6872__132 vssd1 vssd1 vccd1 vccd1 _6872__132/HI _6981_/A sky130_fd_sc_hd__conb_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4770_ _6403_/Q _4778_/B vssd1 vssd1 vccd1 vccd1 _4771_/A sky130_fd_sc_hd__and2_1
XFILLER_119_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ _3757_/A _3605_/B _3722_/C _3765_/A vssd1 vssd1 vccd1 vccd1 _3724_/A sky130_fd_sc_hd__a22o_1
X_6440_ _6795_/CLK _6440_/D vssd1 vssd1 vccd1 vccd1 _6440_/Q sky130_fd_sc_hd__dfxtp_1
X_3652_ _6652_/Q _6651_/Q _6300_/Q _6299_/Q vssd1 vssd1 vccd1 vccd1 _3653_/B sky130_fd_sc_hd__and4_1
X_6371_ _6763_/CLK _6371_/D vssd1 vssd1 vccd1 vccd1 _6371_/Q sky130_fd_sc_hd__dfxtp_1
X_3583_ _6650_/Q _6299_/Q vssd1 vssd1 vccd1 vccd1 _3585_/A sky130_fd_sc_hd__and2_1
X_5322_ _6224_/A _5320_/X _5321_/Y _5775_/B _6624_/Q vssd1 vssd1 vccd1 vccd1 _5499_/B
+ sky130_fd_sc_hd__a2111o_1
X_5253_ _5253_/A vssd1 vssd1 vccd1 vccd1 _6592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5184_ _5191_/A _5184_/B _5184_/C vssd1 vssd1 vccd1 vccd1 _5185_/A sky130_fd_sc_hd__and3_1
X_4204_ _4205_/A _4205_/B _4205_/C vssd1 vssd1 vccd1 vccd1 _4243_/A sky130_fd_sc_hd__o21a_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4135_ _4135_/A _4135_/B _4135_/C vssd1 vssd1 vccd1 vccd1 _4169_/B sky130_fd_sc_hd__nand3_2
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ _4065_/B _4065_/C _4065_/A vssd1 vssd1 vccd1 vccd1 _4066_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4968_ _4968_/A _4968_/B vssd1 vssd1 vccd1 vccd1 _6539_/D sky130_fd_sc_hd__nor2_1
X_4899_ _6518_/Q _4894_/X _4895_/X input45/X vssd1 vssd1 vccd1 vccd1 _6518_/D sky130_fd_sc_hd__a22o_1
X_3919_ _4149_/B _3979_/D _4262_/A _4083_/A vssd1 vssd1 vccd1 vccd1 _3920_/B sky130_fd_sc_hd__a22oi_1
X_6707_ _6789_/CLK _6707_/D vssd1 vssd1 vccd1 vccd1 _6707_/Q sky130_fd_sc_hd__dfxtp_1
X_6638_ _6532_/Q _6638_/D vssd1 vssd1 vccd1 vccd1 _6638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6569_ _6569_/CLK _6569_/D vssd1 vssd1 vccd1 vccd1 _6907_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6856__116 vssd1 vssd1 vccd1 vccd1 _6856__116/HI _6965_/A sky130_fd_sc_hd__conb_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6835__95 vssd1 vssd1 vccd1 vccd1 _6835__95/HI _6944_/A sky130_fd_sc_hd__conb_1
XFILLER_93_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5940_ _6730_/Q _5918_/X _5939_/X _5933_/X vssd1 vssd1 vccd1 vccd1 _6730_/D sky130_fd_sc_hd__o211a_1
XFILLER_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5871_ _5935_/A vssd1 vssd1 vccd1 vccd1 _5871_/X sky130_fd_sc_hd__buf_2
XFILLER_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4822_ _4822_/A vssd1 vssd1 vccd1 vccd1 _6474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4753_ _4753_/A vssd1 vssd1 vccd1 vccd1 _6443_/D sky130_fd_sc_hd__clkbuf_1
X_3704_ _3679_/X _3665_/X _3702_/X _3703_/Y vssd1 vssd1 vccd1 vccd1 _3709_/B sky130_fd_sc_hd__o211ai_1
X_6423_ _6763_/CLK _6423_/D vssd1 vssd1 vccd1 vccd1 _6423_/Q sky130_fd_sc_hd__dfxtp_1
X_4684_ _6349_/Q _4688_/B vssd1 vssd1 vccd1 vccd1 _4685_/A sky130_fd_sc_hd__and2_1
X_3635_ _3592_/X _3631_/X _3634_/Y vssd1 vssd1 vccd1 vccd1 _6340_/D sky130_fd_sc_hd__o21a_1
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6354_ _6763_/CLK _6354_/D vssd1 vssd1 vccd1 vccd1 _6354_/Q sky130_fd_sc_hd__dfxtp_2
X_3566_ _3565_/A _3565_/B _3565_/C vssd1 vssd1 vccd1 vccd1 _3593_/B sky130_fd_sc_hd__a21oi_1
XFILLER_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5305_ _6616_/Q _5305_/B vssd1 vssd1 vccd1 vccd1 _5306_/A sky130_fd_sc_hd__and2_1
X_3497_ _6326_/Q _6530_/Q _3499_/S vssd1 vssd1 vccd1 vccd1 _3498_/A sky130_fd_sc_hd__mux2_1
X_6285_ _6814_/Q _6267_/X _6284_/Y _6275_/X vssd1 vssd1 vccd1 vccd1 _6814_/D sky130_fd_sc_hd__o211a_1
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5236_ _5236_/A _5236_/B _5236_/C vssd1 vssd1 vccd1 vccd1 _5238_/B sky130_fd_sc_hd__and3_1
XFILLER_102_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5167_ _5167_/A vssd1 vssd1 vccd1 vccd1 _6578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5098_ _6812_/Q _5109_/B vssd1 vssd1 vccd1 vccd1 _5098_/X sky130_fd_sc_hd__or2_1
XFILLER_17_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4118_ _4118_/A _4156_/B _4118_/C vssd1 vssd1 vccd1 vccd1 _4160_/A sky130_fd_sc_hd__and3_1
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4049_ _4049_/A _4049_/B vssd1 vssd1 vccd1 vccd1 _4093_/B sky130_fd_sc_hd__or2_1
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3420_ _6299_/Q vssd1 vssd1 vccd1 vccd1 _3762_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3351_ _6644_/Q vssd1 vssd1 vccd1 vccd1 _5406_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3282_ _3286_/A vssd1 vssd1 vccd1 vccd1 _3282_/Y sky130_fd_sc_hd__inv_2
X_6070_ _6070_/A vssd1 vssd1 vccd1 vccd1 _6070_/X sky130_fd_sc_hd__clkbuf_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5021_ _6893_/A _4945_/X _5020_/X _4352_/X vssd1 vssd1 vccd1 vccd1 _6555_/D sky130_fd_sc_hd__o211a_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6972_ _6972_/A _3274_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5923_ _6485_/Q _5931_/B _5943_/C vssd1 vssd1 vccd1 vccd1 _5923_/X sky130_fd_sc_hd__and3_1
X_5854_ _6716_/Q _5850_/X _5853_/X _5838_/X vssd1 vssd1 vccd1 vccd1 _6716_/D sky130_fd_sc_hd__o211a_1
XFILLER_61_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4805_ _4805_/A vssd1 vssd1 vccd1 vccd1 _6466_/D sky130_fd_sc_hd__clkbuf_1
X_5785_ _6623_/Q _5320_/X _5321_/Y _5775_/B _6624_/Q vssd1 vssd1 vccd1 vccd1 _6224_/C
+ sky130_fd_sc_hd__a2111oi_4
X_4736_ _6388_/Q _4744_/B vssd1 vssd1 vccd1 vccd1 _4737_/A sky130_fd_sc_hd__and2_1
X_4667_ _4667_/A vssd1 vssd1 vccd1 vccd1 _6405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6406_ _6789_/CLK _6406_/D vssd1 vssd1 vccd1 vccd1 _6406_/Q sky130_fd_sc_hd__dfxtp_1
X_3618_ _6649_/Q _3758_/B vssd1 vssd1 vccd1 vccd1 _3619_/B sky130_fd_sc_hd__nand2_1
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4598_ _4598_/A _4598_/B vssd1 vssd1 vccd1 vccd1 _4600_/C sky130_fd_sc_hd__xor2_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6337_ _6789_/CLK _6337_/D vssd1 vssd1 vccd1 vccd1 _6337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3549_ _3569_/C _3549_/B vssd1 vssd1 vccd1 vccd1 _3551_/A sky130_fd_sc_hd__xnor2_1
XFILLER_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6268_ _6268_/A vssd1 vssd1 vccd1 vccd1 _6268_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5219_ _6319_/Q _6318_/Q _6317_/Q _6316_/Q vssd1 vssd1 vccd1 vccd1 _5224_/C sky130_fd_sc_hd__or4_1
XFILLER_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6199_ _6789_/Q _6194_/X _6198_/X _6190_/X vssd1 vssd1 vccd1 vccd1 _6789_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5570_ _6467_/Q vssd1 vssd1 vccd1 vccd1 _5570_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4521_ _4557_/A _4542_/B _4520_/X vssd1 vssd1 vccd1 vccd1 _4524_/A sky130_fd_sc_hd__o21bai_1
X_4452_ _4499_/C _4452_/B vssd1 vssd1 vccd1 vccd1 _4453_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3403_ _3578_/B vssd1 vssd1 vccd1 vccd1 _5217_/D sky130_fd_sc_hd__clkbuf_2
X_4383_ _4349_/A _4350_/A _4349_/B vssd1 vssd1 vccd1 vccd1 _4383_/X sky130_fd_sc_hd__a21o_1
XFILLER_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3334_ input27/X input26/X _3334_/C _3334_/D vssd1 vssd1 vccd1 vccd1 _4979_/D sky130_fd_sc_hd__and4bb_1
X_6122_ _6473_/Q _6107_/X _6070_/A _6113_/X _6489_/Q vssd1 vssd1 vccd1 vccd1 _6122_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _5667_/X _5972_/A _6068_/A _6029_/A vssd1 vssd1 vccd1 vccd1 _6053_/X sky130_fd_sc_hd__o31a_1
X_3265_ _3268_/A vssd1 vssd1 vccd1 vccd1 _3265_/Y sky130_fd_sc_hd__inv_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _6551_/Q _5249_/B vssd1 vssd1 vccd1 vccd1 _5005_/A sky130_fd_sc_hd__and2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3196_ _3200_/A vssd1 vssd1 vccd1 vccd1 _3196_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6955_ _6955_/A _3254_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5906_ _5935_/A vssd1 vssd1 vccd1 vccd1 _5906_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5837_ _6487_/Q _5812_/X _5835_/X _5836_/X _5815_/X vssd1 vssd1 vccd1 vccd1 _5837_/X
+ sky130_fd_sc_hd__a221o_1
X_5768_ _6283_/A _5704_/X _5767_/X vssd1 vssd1 vccd1 vccd1 _5768_/X sky130_fd_sc_hd__a21o_1
X_4719_ _4719_/A vssd1 vssd1 vccd1 vccd1 _6428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5699_ _5735_/A vssd1 vssd1 vccd1 vccd1 _5699_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6740_ _6809_/CLK _6740_/D vssd1 vssd1 vccd1 vccd1 _6740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3952_ _3956_/A _3952_/B vssd1 vssd1 vccd1 vccd1 _3953_/C sky130_fd_sc_hd__nand2_1
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6671_ _6795_/CLK _6671_/D vssd1 vssd1 vccd1 vccd1 _6671_/Q sky130_fd_sc_hd__dfxtp_1
X_3883_ _6656_/Q vssd1 vssd1 vccd1 vccd1 _4013_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5622_ _5669_/S vssd1 vssd1 vccd1 vccd1 _5661_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_117_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5553_ _6449_/Q _5603_/B vssd1 vssd1 vccd1 vccd1 _5553_/X sky130_fd_sc_hd__and2_1
X_4504_ _4501_/Y _4502_/X _4466_/Y _4467_/X vssd1 vssd1 vccd1 vccd1 _4566_/B sky130_fd_sc_hd__o211a_1
X_5484_ _5490_/A _5484_/B vssd1 vssd1 vccd1 vccd1 _5485_/A sky130_fd_sc_hd__and2_1
XFILLER_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4435_ _4436_/B _4436_/C _4436_/A vssd1 vssd1 vccd1 vccd1 _4437_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4366_ _4543_/A _4400_/D _4393_/C _4479_/B vssd1 vssd1 vccd1 vccd1 _4366_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3317_ _6499_/Q _3375_/A vssd1 vssd1 vccd1 vccd1 _6499_/D sky130_fd_sc_hd__xor2_1
X_6105_ _6105_/A vssd1 vssd1 vccd1 vccd1 _6759_/D sky130_fd_sc_hd__clkbuf_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _6666_/Q vssd1 vssd1 vccd1 vccd1 _4477_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3249_/A vssd1 vssd1 vccd1 vccd1 _3248_/Y sky130_fd_sc_hd__inv_2
X_6036_ _6489_/Q _6023_/X _6013_/X _6031_/X vssd1 vssd1 vccd1 vccd1 _6036_/X sky130_fd_sc_hd__a31o_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3179_ input1/X vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__clkinv_4
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6938_ _6938_/A _3234_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4220_ _4220_/A _4220_/B _4220_/C _4220_/D vssd1 vssd1 vccd1 vccd1 _4220_/X sky130_fd_sc_hd__or4_2
XFILLER_68_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4151_ _4151_/A _4151_/B vssd1 vssd1 vccd1 vccd1 _4155_/A sky130_fd_sc_hd__nand2_1
X_4082_ _4081_/A _4081_/B _4081_/C vssd1 vssd1 vccd1 vccd1 _4089_/C sky130_fd_sc_hd__a21o_1
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4984_ _4984_/A vssd1 vssd1 vccd1 vccd1 _6544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6723_ _6809_/CLK _6723_/D vssd1 vssd1 vccd1 vccd1 _6723_/Q sky130_fd_sc_hd__dfxtp_1
X_3935_ _3935_/A vssd1 vssd1 vccd1 vccd1 _6361_/D sky130_fd_sc_hd__clkbuf_1
X_6654_ _6763_/CLK _6654_/D vssd1 vssd1 vccd1 vccd1 _6654_/Q sky130_fd_sc_hd__dfxtp_1
X_3866_ _3866_/A vssd1 vssd1 vccd1 vccd1 _6350_/D sky130_fd_sc_hd__clkbuf_1
X_5605_ _5624_/A _5605_/B vssd1 vssd1 vccd1 vccd1 _5605_/X sky130_fd_sc_hd__or2_1
X_6585_ _6586_/CLK _6585_/D vssd1 vssd1 vccd1 vccd1 _6923_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3797_ _3797_/A vssd1 vssd1 vccd1 vccd1 _3797_/Y sky130_fd_sc_hd__inv_2
X_5536_ _6269_/A vssd1 vssd1 vccd1 vccd1 _6286_/B sky130_fd_sc_hd__buf_2
XFILLER_117_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5467_ _5474_/A _5467_/B vssd1 vssd1 vccd1 vccd1 _5468_/A sky130_fd_sc_hd__and2_1
X_4418_ _4418_/A _4418_/B vssd1 vssd1 vccd1 vccd1 _4418_/Y sky130_fd_sc_hd__nor2_1
X_5398_ _6641_/Q _5412_/B vssd1 vssd1 vccd1 vccd1 _5399_/A sky130_fd_sc_hd__and2_1
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4349_ _4349_/A _4349_/B vssd1 vssd1 vccd1 vccd1 _4350_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6019_ _6001_/X _6017_/X _6018_/X vssd1 vssd1 vccd1 vccd1 _6019_/X sky130_fd_sc_hd__a21o_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3720_ _3789_/A _3789_/B _3720_/C _3720_/D vssd1 vssd1 vccd1 vccd1 _3765_/A sky130_fd_sc_hd__nand4_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3651_ _3727_/B _6300_/Q _3720_/C _3727_/A vssd1 vssd1 vccd1 vccd1 _3653_/A sky130_fd_sc_hd__a22oi_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6370_ _6763_/CLK _6370_/D vssd1 vssd1 vccd1 vccd1 _6370_/Q sky130_fd_sc_hd__dfxtp_1
X_3582_ _3727_/A _3727_/B _3645_/B _6297_/Q vssd1 vssd1 vccd1 vccd1 _3585_/C sky130_fd_sc_hd__nand4_1
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5321_ _5406_/A _6644_/Q _6647_/Q _3349_/X vssd1 vssd1 vccd1 vccd1 _5321_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5252_ _6592_/Q _5260_/B vssd1 vssd1 vccd1 vccd1 _5253_/A sky130_fd_sc_hd__and2_1
X_5183_ _5181_/X _5182_/X _5176_/X vssd1 vssd1 vccd1 vccd1 _5184_/C sky130_fd_sc_hd__a21o_1
X_4203_ _4203_/A _4203_/B vssd1 vssd1 vccd1 vccd1 _4205_/C sky130_fd_sc_hd__xor2_1
XFILLER_110_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4134_ _4131_/Y _4132_/X _4098_/B _4098_/Y vssd1 vssd1 vccd1 vccd1 _4135_/C sky130_fd_sc_hd__o211ai_2
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4065_ _4065_/A _4065_/B _4065_/C vssd1 vssd1 vccd1 vccd1 _4065_/Y sky130_fd_sc_hd__nor3_2
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _6539_/Q _4969_/C _4931_/X vssd1 vssd1 vccd1 vccd1 _4968_/B sky130_fd_sc_hd__o21ai_1
XFILLER_51_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4898_ _6517_/Q _4894_/X _4895_/X input44/X vssd1 vssd1 vccd1 vccd1 _6517_/D sky130_fd_sc_hd__a22o_1
X_6706_ _6789_/CLK _6706_/D vssd1 vssd1 vccd1 vccd1 _6706_/Q sky130_fd_sc_hd__dfxtp_1
X_3918_ _4149_/B _6658_/Q _4039_/C _4039_/D vssd1 vssd1 vccd1 vccd1 _3957_/C sky130_fd_sc_hd__and4_1
X_6637_ _6799_/CLK _6637_/D vssd1 vssd1 vccd1 vccd1 _6637_/Q sky130_fd_sc_hd__dfxtp_1
X_3849_ _3849_/A _3879_/A vssd1 vssd1 vccd1 vccd1 _3850_/C sky130_fd_sc_hd__nand2_1
X_6568_ _6569_/CLK _6568_/D vssd1 vssd1 vccd1 vccd1 _6906_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5519_ _6031_/A vssd1 vssd1 vccd1 vccd1 _5519_/X sky130_fd_sc_hd__buf_2
X_6499_ _6554_/CLK _6499_/D hold3/A vssd1 vssd1 vccd1 vccd1 _6499_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _5870_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__or2_2
XFILLER_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4821_ _6426_/Q _4823_/B vssd1 vssd1 vccd1 vccd1 _4822_/A sky130_fd_sc_hd__and2_1
XFILLER_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ _6395_/Q _4756_/B vssd1 vssd1 vccd1 vccd1 _4753_/A sky130_fd_sc_hd__and2_1
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3703_ _3703_/A _3703_/B _3703_/C vssd1 vssd1 vccd1 vccd1 _3703_/Y sky130_fd_sc_hd__nand3_2
X_4683_ _4683_/A vssd1 vssd1 vccd1 vccd1 _6412_/D sky130_fd_sc_hd__clkbuf_1
X_3634_ _3592_/X _3631_/X _3633_/X vssd1 vssd1 vccd1 vccd1 _3634_/Y sky130_fd_sc_hd__a21oi_1
X_6422_ _6763_/CLK _6422_/D vssd1 vssd1 vccd1 vccd1 _6422_/Q sky130_fd_sc_hd__dfxtp_1
X_6353_ _6763_/CLK _6353_/D vssd1 vssd1 vccd1 vccd1 _6353_/Q sky130_fd_sc_hd__dfxtp_1
X_3565_ _3565_/A _3565_/B _3565_/C vssd1 vssd1 vccd1 vccd1 _3567_/B sky130_fd_sc_hd__and3_1
X_5304_ _5304_/A vssd1 vssd1 vccd1 vccd1 _6615_/D sky130_fd_sc_hd__clkbuf_1
X_3496_ _3496_/A vssd1 vssd1 vccd1 vccd1 _6325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6284_ _6268_/X _6283_/Y _6267_/A vssd1 vssd1 vccd1 vccd1 _6284_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5235_ _5414_/C _5235_/B _5235_/C vssd1 vssd1 vccd1 vccd1 _5236_/C sky130_fd_sc_hd__nor3_1
XFILLER_102_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5166_ _5191_/A _5166_/B _5166_/C vssd1 vssd1 vccd1 vccd1 _5167_/A sky130_fd_sc_hd__and3_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5097_ _5108_/A _5097_/B vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__or2_1
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4117_ _4079_/A _4079_/B _4079_/C vssd1 vssd1 vccd1 vccd1 _4118_/C sky130_fd_sc_hd__a21bo_1
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6879__139 vssd1 vssd1 vccd1 vccd1 _6879__139/HI _6988_/A sky130_fd_sc_hd__conb_1
XFILLER_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4048_ _4121_/A _4121_/B _4153_/C _6354_/Q vssd1 vssd1 vccd1 vccd1 _4049_/B sky130_fd_sc_hd__and4_1
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _5999_/A vssd1 vssd1 vccd1 vccd1 _5999_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3350_ _6645_/Q vssd1 vssd1 vccd1 vccd1 _5406_/A sky130_fd_sc_hd__buf_2
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3281_/A vssd1 vssd1 vccd1 vccd1 _3286_/A sky130_fd_sc_hd__buf_12
X_5020_ _5011_/X _5016_/X _5019_/X vssd1 vssd1 vccd1 vccd1 _5020_/X sky130_fd_sc_hd__a21o_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6971_ _6971_/A _3273_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
XFILLER_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5922_ _5922_/A vssd1 vssd1 vccd1 vccd1 _5943_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5853_ _6490_/Q _5840_/X _5852_/X _5836_/X _5843_/X vssd1 vssd1 vccd1 vccd1 _5853_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4804_ _6418_/Q _4812_/B vssd1 vssd1 vccd1 vccd1 _4805_/A sky130_fd_sc_hd__and2_1
X_5784_ _5506_/X _5780_/X _5860_/S vssd1 vssd1 vccd1 vccd1 _5784_/X sky130_fd_sc_hd__mux2_1
X_4735_ _4735_/A vssd1 vssd1 vccd1 vccd1 _4744_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4666_ _6341_/Q _4666_/B vssd1 vssd1 vccd1 vccd1 _4667_/A sky130_fd_sc_hd__and2_1
X_4597_ _4597_/A _4597_/B vssd1 vssd1 vccd1 vccd1 _4598_/B sky130_fd_sc_hd__nand2_1
X_3617_ _3585_/A _3585_/B _3585_/C vssd1 vssd1 vccd1 vccd1 _3638_/C sky130_fd_sc_hd__a21bo_1
X_6405_ _6789_/CLK _6405_/D vssd1 vssd1 vccd1 vccd1 _6405_/Q sky130_fd_sc_hd__dfxtp_1
X_3548_ _4385_/A vssd1 vssd1 vccd1 vccd1 _6067_/A sky130_fd_sc_hd__buf_4
X_6336_ _6763_/CLK _6336_/D vssd1 vssd1 vccd1 vccd1 _6336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6267_ _6267_/A vssd1 vssd1 vccd1 vccd1 _6267_/X sky130_fd_sc_hd__clkbuf_2
X_3479_ _3479_/A vssd1 vssd1 vccd1 vccd1 _6317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5218_ _5218_/A _5218_/B _5218_/C vssd1 vssd1 vccd1 vccd1 _5224_/B sky130_fd_sc_hd__or3_1
X_6198_ _6250_/A _6205_/B vssd1 vssd1 vccd1 vccd1 _6198_/X sky130_fd_sc_hd__or2_1
X_5149_ _6914_/A _5149_/B vssd1 vssd1 vccd1 vccd1 _5153_/B sky130_fd_sc_hd__or2_1
XFILLER_84_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4520_ _4541_/A _4541_/B vssd1 vssd1 vccd1 vccd1 _4520_/X sky130_fd_sc_hd__xor2_1
X_4451_ _4451_/A _4579_/B vssd1 vssd1 vccd1 vccd1 _4452_/B sky130_fd_sc_hd__nand2_1
X_3402_ _6296_/Q vssd1 vssd1 vccd1 vccd1 _3578_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4382_ _4382_/A _4382_/B vssd1 vssd1 vccd1 vccd1 _4382_/X sky130_fd_sc_hd__or2_1
X_6121_ _6121_/A vssd1 vssd1 vccd1 vccd1 _6762_/D sky130_fd_sc_hd__clkbuf_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3333_ _3333_/A _3333_/B _3333_/C _3333_/D vssd1 vssd1 vccd1 vccd1 _4979_/C sky130_fd_sc_hd__nor4_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6052_ _6750_/Q _5523_/X _6050_/X _6051_/X vssd1 vssd1 vccd1 vccd1 _6750_/D sky130_fd_sc_hd__o211a_1
X_3264_ _3268_/A vssd1 vssd1 vccd1 vccd1 _3264_/Y sky130_fd_sc_hd__inv_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5003_ _5879_/A _5003_/B vssd1 vssd1 vccd1 vccd1 _6550_/D sky130_fd_sc_hd__nor2_1
XFILLER_100_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _3219_/A vssd1 vssd1 vccd1 vccd1 _3200_/A sky130_fd_sc_hd__buf_4
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6954_ _6954_/A _3253_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5905_ _6724_/Q _5888_/X _5903_/X _5904_/X vssd1 vssd1 vccd1 vccd1 _6724_/D sky130_fd_sc_hd__o211a_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5836_ _5836_/A vssd1 vssd1 vccd1 vccd1 _5836_/X sky130_fd_sc_hd__clkbuf_2
X_5767_ _5915_/A vssd1 vssd1 vccd1 vccd1 _5767_/X sky130_fd_sc_hd__clkbuf_2
X_4718_ _6372_/Q _4722_/B vssd1 vssd1 vccd1 vccd1 _4719_/A sky130_fd_sc_hd__and2_1
X_5698_ _5721_/S vssd1 vssd1 vccd1 vccd1 _5698_/X sky130_fd_sc_hd__clkbuf_2
X_4649_ _4637_/A _4637_/B _4648_/X _4644_/A vssd1 vssd1 vccd1 vccd1 _4649_/X sky130_fd_sc_hd__a31o_1
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6319_ _6523_/CLK _6319_/D vssd1 vssd1 vccd1 vccd1 _6319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3951_ _3951_/A _3951_/B vssd1 vssd1 vccd1 vccd1 _3952_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6670_ _6795_/CLK _6670_/D vssd1 vssd1 vccd1 vccd1 _6670_/Q sky130_fd_sc_hd__dfxtp_1
X_3882_ _3882_/A vssd1 vssd1 vccd1 vccd1 _6357_/D sky130_fd_sc_hd__clkbuf_1
X_5621_ _6456_/Q _5660_/B vssd1 vssd1 vccd1 vccd1 _5621_/X sky130_fd_sc_hd__and2_2
XFILLER_31_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5552_ _6465_/Q vssd1 vssd1 vccd1 vccd1 _5552_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4503_ _4466_/Y _4467_/X _4501_/Y _4502_/X vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__a211oi_4
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5483_ _6315_/Q _4545_/B _5483_/S vssd1 vssd1 vccd1 vccd1 _5484_/B sky130_fd_sc_hd__mux2_1
X_4434_ _6669_/Q _4510_/C vssd1 vssd1 vccd1 vccd1 _4436_/A sky130_fd_sc_hd__and2_1
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4365_ _4517_/A vssd1 vssd1 vccd1 vccd1 _4543_/A sky130_fd_sc_hd__clkbuf_2
X_3316_ _6498_/Q _6497_/Q _3373_/B vssd1 vssd1 vccd1 vccd1 _3375_/A sky130_fd_sc_hd__and3_1
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _6110_/A _6104_/B vssd1 vssd1 vccd1 vccd1 _6105_/A sky130_fd_sc_hd__and2_1
X_4296_ _4296_/A _4407_/A _4296_/C _4333_/B vssd1 vssd1 vccd1 vccd1 _4296_/X sky130_fd_sc_hd__and4_1
X_6035_ _6747_/Q _5630_/X _6044_/S vssd1 vssd1 vccd1 vccd1 _6035_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3249_/A vssd1 vssd1 vccd1 vccd1 _3247_/Y sky130_fd_sc_hd__inv_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6937_ _6937_/A _3233_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5819_ _6710_/Q _5584_/X _5841_/S vssd1 vssd1 vccd1 vccd1 _5819_/X sky130_fd_sc_hd__mux2_1
X_6799_ _6799_/CLK _6799_/D vssd1 vssd1 vccd1 vccd1 _6799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4150_ _4150_/A _4192_/A vssd1 vssd1 vccd1 vccd1 _4188_/A sky130_fd_sc_hd__or2_1
XFILLER_95_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4081_ _4081_/A _4081_/B _4081_/C vssd1 vssd1 vccd1 vccd1 _4089_/B sky130_fd_sc_hd__nand3_1
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4983_ _4986_/B _5239_/B _4983_/C vssd1 vssd1 vccd1 vccd1 _4984_/A sky130_fd_sc_hd__and3b_1
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6722_ _6809_/CLK _6722_/D vssd1 vssd1 vccd1 vccd1 _6722_/Q sky130_fd_sc_hd__dfxtp_1
X_3934_ _4325_/A _3934_/B _3953_/B vssd1 vssd1 vccd1 vccd1 _3935_/A sky130_fd_sc_hd__and3_1
X_6653_ _6763_/CLK _6653_/D vssd1 vssd1 vccd1 vccd1 _6653_/Q sky130_fd_sc_hd__dfxtp_1
X_3865_ _3865_/A _6275_/A vssd1 vssd1 vccd1 vccd1 _3866_/A sky130_fd_sc_hd__and2_1
X_5604_ _6680_/Q _5603_/X _5612_/S vssd1 vssd1 vccd1 vccd1 _5605_/B sky130_fd_sc_hd__mux2_1
X_6584_ _6584_/CLK _6584_/D vssd1 vssd1 vccd1 vccd1 _6922_/A sky130_fd_sc_hd__dfxtp_1
X_3796_ _3796_/A _3796_/B vssd1 vssd1 vccd1 vccd1 _3820_/A sky130_fd_sc_hd__xnor2_2
X_5535_ _5535_/A vssd1 vssd1 vccd1 vccd1 _6269_/A sky130_fd_sc_hd__buf_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5466_ _6310_/Q _4241_/A _5466_/S vssd1 vssd1 vccd1 vccd1 _5467_/B sky130_fd_sc_hd__mux2_1
X_4417_ _4416_/B _4416_/C _4416_/A vssd1 vssd1 vccd1 vccd1 _4420_/B sky130_fd_sc_hd__a21o_1
X_5397_ _5397_/A vssd1 vssd1 vccd1 vccd1 _6640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4348_ _4348_/A _4348_/B vssd1 vssd1 vccd1 vccd1 _4349_/B sky130_fd_sc_hd__or2_1
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4279_ _4449_/A vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6018_ _6486_/Q _5996_/X _6013_/X _6003_/X vssd1 vssd1 vccd1 vccd1 _6018_/X sky130_fd_sc_hd__a31o_1
XFILLER_100_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3650_ _3650_/A _3758_/B vssd1 vssd1 vccd1 vccd1 _3698_/A sky130_fd_sc_hd__nand2_1
X_3581_ _6298_/Q vssd1 vssd1 vccd1 vccd1 _3645_/B sky130_fd_sc_hd__clkbuf_2
X_5320_ _6622_/Q _6621_/Q _5880_/B vssd1 vssd1 vccd1 vccd1 _5320_/X sky130_fd_sc_hd__or3_1
X_5251_ _5273_/A vssd1 vssd1 vccd1 vccd1 _5260_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4202_ _4202_/A _4230_/D vssd1 vssd1 vccd1 vccd1 _4203_/B sky130_fd_sc_hd__nand2_1
XFILLER_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5182_ _6698_/Q _6730_/Q _6762_/Q _6794_/Q _5157_/X _5169_/X vssd1 vssd1 vccd1 vccd1
+ _5182_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4133_ _4098_/B _4098_/Y _4131_/Y _4132_/X vssd1 vssd1 vccd1 vccd1 _4135_/B sky130_fd_sc_hd__a211o_1
XFILLER_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ _4061_/Y _4062_/X _4019_/B _4035_/Y vssd1 vssd1 vccd1 vccd1 _4065_/C sky130_fd_sc_hd__o211a_1
XFILLER_95_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4966_ _6539_/Q _4969_/C vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__and2_1
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6705_ _6789_/CLK _6705_/D vssd1 vssd1 vccd1 vccd1 _6705_/Q sky130_fd_sc_hd__dfxtp_1
X_4897_ _6516_/Q _4894_/X _4895_/X input43/X vssd1 vssd1 vccd1 vccd1 _6516_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3917_ _3944_/B vssd1 vssd1 vccd1 vccd1 _4149_/B sky130_fd_sc_hd__clkbuf_2
X_6636_ _6799_/CLK _6636_/D vssd1 vssd1 vccd1 vccd1 _6636_/Q sky130_fd_sc_hd__dfxtp_1
X_3848_ _3843_/A _3847_/Y _3843_/B vssd1 vssd1 vccd1 vccd1 _3848_/Y sky130_fd_sc_hd__o21ai_1
X_6567_ _6569_/CLK _6567_/D vssd1 vssd1 vccd1 vccd1 _6905_/A sky130_fd_sc_hd__dfxtp_1
X_3779_ _3718_/X _3745_/Y _3778_/C vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5518_ _5518_/A vssd1 vssd1 vccd1 vccd1 _6031_/A sky130_fd_sc_hd__buf_2
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6523_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6498_ _6554_/CLK _6498_/D hold3/A vssd1 vssd1 vccd1 vccd1 _6498_/Q sky130_fd_sc_hd__dfrtp_1
X_5449_ _5456_/A _5449_/B vssd1 vssd1 vccd1 vccd1 _5450_/A sky130_fd_sc_hd__and2_1
XFILLER_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4820_ _4820_/A vssd1 vssd1 vccd1 vccd1 _6473_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4751_/A vssd1 vssd1 vccd1 vccd1 _6442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3702_ _3703_/B _3703_/C _3703_/A vssd1 vssd1 vccd1 vccd1 _3702_/X sky130_fd_sc_hd__a21o_1
X_4682_ _6348_/Q _4688_/B vssd1 vssd1 vccd1 vccd1 _4683_/A sky130_fd_sc_hd__and2_1
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3633_ _3636_/A vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__buf_4
X_6421_ _6763_/CLK _6421_/D vssd1 vssd1 vccd1 vccd1 _6421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6352_ _6763_/CLK _6352_/D vssd1 vssd1 vccd1 vccd1 _6352_/Q sky130_fd_sc_hd__dfxtp_1
X_3564_ _3568_/A _3564_/B vssd1 vssd1 vccd1 vccd1 _3565_/C sky130_fd_sc_hd__nand2_1
X_5303_ _6615_/Q _5305_/B vssd1 vssd1 vccd1 vccd1 _5304_/A sky130_fd_sc_hd__and2_1
X_3495_ _6325_/Q _6529_/Q _3495_/S vssd1 vssd1 vccd1 vccd1 _3496_/A sky130_fd_sc_hd__mux2_1
X_6283_ _6283_/A _6283_/B vssd1 vssd1 vccd1 vccd1 _6283_/Y sky130_fd_sc_hd__nand2_1
X_5234_ _6619_/Q _6618_/Q _6617_/Q _6616_/Q vssd1 vssd1 vccd1 vccd1 _5235_/C sky130_fd_sc_hd__or4_1
XFILLER_102_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5165_ _5150_/X _5164_/X _5145_/X vssd1 vssd1 vccd1 vccd1 _5166_/C sky130_fd_sc_hd__a21o_1
XFILLER_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4116_ _4151_/A _4116_/B _4116_/C _4156_/A vssd1 vssd1 vccd1 vccd1 _4156_/B sky130_fd_sc_hd__nand4_2
X_5096_ _6684_/Q _6716_/Q _6748_/Q _6780_/Q _5083_/X _4949_/A vssd1 vssd1 vccd1 vccd1
+ _5097_/B sky130_fd_sc_hd__mux4_1
XFILLER_56_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6826__86 vssd1 vssd1 vccd1 vccd1 _6826__86/HI _6935_/A sky130_fd_sc_hd__conb_1
XFILLER_17_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4047_ _4147_/A _3998_/D _4180_/C _4085_/B vssd1 vssd1 vccd1 vccd1 _4049_/A sky130_fd_sc_hd__a22oi_1
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5969_/X _5995_/X _5997_/X vssd1 vssd1 vccd1 vccd1 _5998_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4949_ _4949_/A vssd1 vssd1 vccd1 vccd1 _4950_/A sky130_fd_sc_hd__clkbuf_4
X_6619_ _6667_/CLK _6619_/D vssd1 vssd1 vccd1 vccd1 _6619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6862__122 vssd1 vssd1 vccd1 vccd1 _6862__122/HI _6971_/A sky130_fd_sc_hd__conb_1
XFILLER_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3280_ _3280_/A vssd1 vssd1 vccd1 vccd1 _3280_/Y sky130_fd_sc_hd__inv_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6970_ _6970_/A _3272_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
XFILLER_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _5593_/X _5919_/X _5920_/X _5912_/X _6727_/Q vssd1 vssd1 vccd1 vccd1 _5921_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5852_ _5642_/X _5851_/X _5860_/S vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__mux2_1
X_5783_ _5866_/S vssd1 vssd1 vccd1 vccd1 _5860_/S sky130_fd_sc_hd__buf_2
X_4803_ _4847_/A vssd1 vssd1 vccd1 vccd1 _4812_/B sky130_fd_sc_hd__clkbuf_1
X_4734_ _4734_/A vssd1 vssd1 vccd1 vccd1 _6435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4665_ _4665_/A vssd1 vssd1 vccd1 vccd1 _6404_/D sky130_fd_sc_hd__clkbuf_1
X_4596_ _4596_/A _4596_/B vssd1 vssd1 vccd1 vccd1 _4598_/A sky130_fd_sc_hd__nand2_1
X_3616_ _3616_/A _3755_/D vssd1 vssd1 vccd1 vccd1 _3620_/A sky130_fd_sc_hd__nand2_1
X_6404_ _6789_/CLK _6404_/D vssd1 vssd1 vccd1 vccd1 _6404_/Q sky130_fd_sc_hd__dfxtp_1
X_3547_ _3632_/A vssd1 vssd1 vccd1 vccd1 _4385_/A sky130_fd_sc_hd__buf_2
X_6335_ _6763_/CLK _6335_/D vssd1 vssd1 vccd1 vccd1 _6335_/Q sky130_fd_sc_hd__dfxtp_1
X_6846__106 vssd1 vssd1 vccd1 vccd1 _6846__106/HI _6955_/A sky130_fd_sc_hd__conb_1
X_3478_ _6317_/Q _6521_/Q _3484_/S vssd1 vssd1 vccd1 vccd1 _3479_/A sky130_fd_sc_hd__mux2_1
X_6266_ _6809_/Q _6247_/X _6265_/Y _6255_/X vssd1 vssd1 vccd1 vccd1 _6809_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5217_ _5217_/A _5217_/B _5217_/C _5217_/D vssd1 vssd1 vccd1 vccd1 _5218_/C sky130_fd_sc_hd__or4_2
X_6197_ _6788_/Q _6194_/X _6196_/X _6190_/X vssd1 vssd1 vccd1 vccd1 _6788_/D sky130_fd_sc_hd__o211a_1
X_5148_ _5148_/A vssd1 vssd1 vccd1 vccd1 _6575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _5047_/X _5077_/X _5078_/X _5055_/X vssd1 vssd1 vccd1 vccd1 _5079_/X sky130_fd_sc_hd__a31o_2
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _4450_/A _4450_/B vssd1 vssd1 vccd1 vccd1 _4499_/C sky130_fd_sc_hd__nand2_1
XFILLER_109_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3401_ _6295_/Q _3396_/X _3400_/Y vssd1 vssd1 vccd1 vccd1 _6295_/D sky130_fd_sc_hd__o21a_1
X_4381_ _4381_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4382_/B sky130_fd_sc_hd__and2_1
XFILLER_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3332_ _3332_/A _3332_/B vssd1 vssd1 vccd1 vccd1 _4979_/B sky130_fd_sc_hd__nor2_1
X_6120_ _6132_/A _6120_/B vssd1 vssd1 vccd1 vccd1 _6121_/A sky130_fd_sc_hd__and2_1
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3281_/A vssd1 vssd1 vccd1 vccd1 _3268_/A sky130_fd_sc_hd__buf_12
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6051_ _6178_/A vssd1 vssd1 vccd1 vccd1 _6051_/X sky130_fd_sc_hd__clkbuf_4
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _6549_/Q _4998_/B _6550_/Q vssd1 vssd1 vccd1 vccd1 _5003_/B sky130_fd_sc_hd__a21oi_1
X_3194_ input1/X vssd1 vssd1 vccd1 vccd1 _3219_/A sky130_fd_sc_hd__clkbuf_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6953_ _6953_/A _3252_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
X_5904_ _5999_/A vssd1 vssd1 vccd1 vccd1 _5904_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5835_ _5610_/X _5834_/X _5842_/S vssd1 vssd1 vccd1 vccd1 _5835_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5766_ _5659_/X _5698_/X _5735_/A _5765_/X vssd1 vssd1 vccd1 vccd1 _5766_/X sky130_fd_sc_hd__o211a_1
XFILLER_10_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4717_ _4717_/A vssd1 vssd1 vccd1 vccd1 _6427_/D sky130_fd_sc_hd__clkbuf_1
X_5697_ _6689_/Q _3357_/X _5696_/X _5690_/X vssd1 vssd1 vccd1 vccd1 _6689_/D sky130_fd_sc_hd__o211a_1
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4648_ _4636_/A _4636_/B _4640_/B vssd1 vssd1 vccd1 vccd1 _4648_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4579_ _4597_/A _4579_/B _4579_/C vssd1 vssd1 vccd1 vccd1 _4600_/B sky130_fd_sc_hd__and3_1
X_6318_ _6523_/CLK _6318_/D vssd1 vssd1 vccd1 vccd1 _6318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6249_ _6249_/A vssd1 vssd1 vccd1 vccd1 _6263_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6586_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_67_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3950_ _3951_/A _3951_/B vssd1 vssd1 vccd1 vccd1 _3956_/A sky130_fd_sc_hd__or2_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3881_ _3881_/A _4257_/B vssd1 vssd1 vccd1 vccd1 _3882_/A sky130_fd_sc_hd__and2_1
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5620_ _5620_/A vssd1 vssd1 vccd1 vccd1 _5620_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5551_ _5650_/A vssd1 vssd1 vccd1 vccd1 _5551_/X sky130_fd_sc_hd__clkbuf_2
X_4502_ _4502_/A _4502_/B _4502_/C vssd1 vssd1 vccd1 vccd1 _4502_/X sky130_fd_sc_hd__and3_1
XFILLER_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5482_ _5482_/A vssd1 vssd1 vccd1 vccd1 _6666_/D sky130_fd_sc_hd__clkbuf_1
X_4433_ _4576_/A _4510_/B _4433_/C _4433_/D vssd1 vssd1 vccd1 vccd1 _4436_/C sky130_fd_sc_hd__nand4_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4364_ _6668_/Q vssd1 vssd1 vccd1 vccd1 _4517_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3315_ _6496_/Q _6495_/Q _3370_/B vssd1 vssd1 vccd1 vccd1 _3373_/B sky130_fd_sc_hd__and3_1
XFILLER_112_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4295_ _4393_/C vssd1 vssd1 vccd1 vccd1 _4333_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6103_ _6759_/Q _6080_/X _6101_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6104_/B sky130_fd_sc_hd__a22o_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3249_/A vssd1 vssd1 vccd1 vccd1 _3246_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6034_ _6746_/Q _6011_/X _6033_/X _6027_/X vssd1 vssd1 vccd1 vccd1 _6746_/D sky130_fd_sc_hd__o211a_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6936_ _6936_/A _3231_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6798_ _6799_/CLK _6798_/D vssd1 vssd1 vccd1 vccd1 _6798_/Q sky130_fd_sc_hd__dfxtp_1
X_5818_ _5865_/S vssd1 vssd1 vccd1 vccd1 _5841_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_50_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5749_ _6270_/A _5704_/X _5705_/X vssd1 vssd1 vccd1 vccd1 _5749_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4080_ _4042_/A _4042_/B _4042_/C vssd1 vssd1 vccd1 vccd1 _4081_/C sky130_fd_sc_hd__a21bo_1
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4982_ _6544_/Q _4982_/B vssd1 vssd1 vccd1 vccd1 _4983_/C sky130_fd_sc_hd__or2_1
X_6721_ _6809_/CLK _6721_/D vssd1 vssd1 vccd1 vccd1 _6721_/Q sky130_fd_sc_hd__dfxtp_1
X_3933_ _3933_/A _3933_/B vssd1 vssd1 vccd1 vccd1 _3953_/B sky130_fd_sc_hd__or2_1
X_3864_ _5193_/A vssd1 vssd1 vccd1 vccd1 _6275_/A sky130_fd_sc_hd__buf_6
X_6652_ _6763_/CLK _6652_/D vssd1 vssd1 vccd1 vccd1 _6652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5603_ _6454_/Q _5603_/B vssd1 vssd1 vccd1 vccd1 _5603_/X sky130_fd_sc_hd__and2_2
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6583_ _6586_/CLK _6583_/D vssd1 vssd1 vccd1 vccd1 _6921_/A sky130_fd_sc_hd__dfxtp_4
X_3795_ _3815_/B _3795_/B vssd1 vssd1 vccd1 vccd1 _3796_/B sky130_fd_sc_hd__xnor2_2
XFILLER_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5534_ _5638_/A vssd1 vssd1 vccd1 vccd1 _5534_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5465_ _5465_/A vssd1 vssd1 vccd1 vccd1 _6661_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4416_ _4416_/A _4416_/B _4416_/C vssd1 vssd1 vccd1 vccd1 _4420_/A sky130_fd_sc_hd__nand3_2
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5396_ _6640_/Q _5396_/B vssd1 vssd1 vccd1 vccd1 _5397_/A sky130_fd_sc_hd__and2_1
XFILLER_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4347_ _4347_/A _4347_/B vssd1 vssd1 vccd1 vccd1 _4348_/B sky130_fd_sc_hd__nor2_1
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4278_ _4407_/A vssd1 vssd1 vccd1 vccd1 _4449_/A sky130_fd_sc_hd__clkbuf_2
X_3229_ _3231_/A vssd1 vssd1 vccd1 vccd1 _3229_/Y sky130_fd_sc_hd__inv_2
X_6017_ _6744_/Q _5602_/X _6017_/S vssd1 vssd1 vccd1 vccd1 _6017_/X sky130_fd_sc_hd__mux2_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6919_ _6919_/A _3211_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__ebufn_8
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3580_ _6652_/Q vssd1 vssd1 vccd1 vccd1 _3727_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5250_ _5250_/A vssd1 vssd1 vccd1 vccd1 _6591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4201_ _4201_/A _4201_/B vssd1 vssd1 vccd1 vccd1 _4203_/A sky130_fd_sc_hd__nand2_1
X_5181_ _5181_/A vssd1 vssd1 vccd1 vccd1 _5181_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4132_ _4144_/A _4144_/B _4144_/C vssd1 vssd1 vccd1 vccd1 _4132_/X sky130_fd_sc_hd__and3_1
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4063_ _4019_/B _4035_/Y _4061_/Y _4062_/X vssd1 vssd1 vccd1 vccd1 _4065_/B sky130_fd_sc_hd__a211oi_4
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4965_ _4965_/A vssd1 vssd1 vccd1 vccd1 _6538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3916_ _6659_/Q vssd1 vssd1 vccd1 vccd1 _3944_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6704_ _6809_/CLK _6704_/D vssd1 vssd1 vccd1 vccd1 _6704_/Q sky130_fd_sc_hd__dfxtp_1
X_4896_ _6515_/Q _4894_/X _4895_/X input42/X vssd1 vssd1 vccd1 vccd1 _6515_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6635_ _6532_/Q _6635_/D vssd1 vssd1 vccd1 vccd1 _6635_/Q sky130_fd_sc_hd__dfxtp_1
X_3847_ _3847_/A vssd1 vssd1 vccd1 vccd1 _3847_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6566_ _6569_/CLK _6566_/D vssd1 vssd1 vccd1 vccd1 _6904_/A sky130_fd_sc_hd__dfxtp_1
X_3778_ _3778_/A _3778_/B _3778_/C _3745_/Y vssd1 vssd1 vccd1 vccd1 _3828_/C sky130_fd_sc_hd__or4b_1
X_5517_ _6040_/A vssd1 vssd1 vccd1 vccd1 _6056_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6497_ _6554_/CLK _6497_/D hold3/A vssd1 vssd1 vccd1 vccd1 _6497_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5448_ _6305_/Q _4103_/A _5448_/S vssd1 vssd1 vccd1 vccd1 _5449_/B sky130_fd_sc_hd__mux2_1
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5379_ _6102_/A vssd1 vssd1 vccd1 vccd1 _5650_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _6394_/Q _4756_/B vssd1 vssd1 vccd1 vccd1 _4751_/A sky130_fd_sc_hd__and2_1
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3701_ _3741_/A _3701_/B vssd1 vssd1 vccd1 vccd1 _3703_/A sky130_fd_sc_hd__nor2_1
X_4681_ _4681_/A vssd1 vssd1 vccd1 vccd1 _6411_/D sky130_fd_sc_hd__clkbuf_1
X_3632_ _3632_/A vssd1 vssd1 vccd1 vccd1 _3636_/A sky130_fd_sc_hd__buf_4
X_6420_ _6763_/CLK _6420_/D vssd1 vssd1 vccd1 vccd1 _6420_/Q sky130_fd_sc_hd__dfxtp_1
X_6351_ _6763_/CLK _6351_/D vssd1 vssd1 vccd1 vccd1 _6351_/Q sky130_fd_sc_hd__dfxtp_1
X_5302_ _5302_/A vssd1 vssd1 vccd1 vccd1 _6614_/D sky130_fd_sc_hd__clkbuf_1
X_3563_ _3563_/A _3563_/B vssd1 vssd1 vccd1 vccd1 _3564_/B sky130_fd_sc_hd__nand2_1
X_3494_ _3494_/A vssd1 vssd1 vccd1 vccd1 _6324_/D sky130_fd_sc_hd__clkbuf_1
X_6282_ _6813_/Q _6267_/X _6281_/Y _6275_/X vssd1 vssd1 vccd1 vccd1 _6813_/D sky130_fd_sc_hd__o211a_1
X_5233_ _6615_/Q _6604_/Q _6589_/Q _6328_/Q vssd1 vssd1 vccd1 vccd1 _5235_/B sky130_fd_sc_hd__or4b_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5164_ _6695_/Q _6727_/Q _6759_/Q _6791_/Q _5157_/X _5138_/X vssd1 vssd1 vccd1 vccd1
+ _5164_/X sky130_fd_sc_hd__mux4_2
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4115_ _6661_/Q _4180_/C _4116_/C _4156_/A vssd1 vssd1 vccd1 vccd1 _4118_/A sky130_fd_sc_hd__a22o_1
X_5095_ _6904_/A _5075_/X _5094_/X _5068_/X vssd1 vssd1 vccd1 vccd1 _6566_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4046_ _6354_/Q vssd1 vssd1 vccd1 vccd1 _4180_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_17_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _6482_/Q _5996_/X _5986_/X _5976_/X vssd1 vssd1 vccd1 vccd1 _5997_/X sky130_fd_sc_hd__a31o_1
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4948_ _6534_/Q vssd1 vssd1 vccd1 vccd1 _4949_/A sky130_fd_sc_hd__clkbuf_2
X_4879_ _4929_/S vssd1 vssd1 vccd1 vccd1 _4910_/S sky130_fd_sc_hd__buf_4
X_6618_ _6667_/CLK _6618_/D vssd1 vssd1 vccd1 vccd1 _6618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6549_ _6551_/CLK _6549_/D vssd1 vssd1 vccd1 vccd1 _6549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5920_ _5920_/A vssd1 vssd1 vccd1 vccd1 _5920_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5851_ _6716_/Q _5643_/X _5859_/S vssd1 vssd1 vccd1 vccd1 _5851_/X sky130_fd_sc_hd__mux2_1
X_5782_ _5882_/A _5872_/A _5872_/B vssd1 vssd1 vccd1 vccd1 _5866_/S sky130_fd_sc_hd__or3_4
X_4802_ _5284_/A vssd1 vssd1 vccd1 vccd1 _4847_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4733_ _6387_/Q _4733_/B vssd1 vssd1 vccd1 vccd1 _4734_/A sky130_fd_sc_hd__and2_1
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4664_ _6340_/Q _4666_/B vssd1 vssd1 vccd1 vccd1 _4665_/A sky130_fd_sc_hd__and2_1
X_6403_ _6789_/CLK _6403_/D vssd1 vssd1 vccd1 vccd1 _6403_/Q sky130_fd_sc_hd__dfxtp_1
X_4595_ _4622_/A _4623_/A _4595_/C _4595_/D vssd1 vssd1 vccd1 vccd1 _4596_/B sky130_fd_sc_hd__nand4_1
X_3615_ _3614_/B _3614_/C _3614_/A vssd1 vssd1 vccd1 vccd1 _3622_/C sky130_fd_sc_hd__a21o_1
X_6885__145 vssd1 vssd1 vccd1 vccd1 _6885__145/HI _6994_/A sky130_fd_sc_hd__conb_1
XFILLER_115_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3546_ _3546_/A vssd1 vssd1 vccd1 vccd1 _6337_/D sky130_fd_sc_hd__clkbuf_1
X_6334_ _6763_/CLK _6334_/D vssd1 vssd1 vccd1 vccd1 _6334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6265_ _6248_/X _6263_/Y _6264_/X vssd1 vssd1 vccd1 vccd1 _6265_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_103_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3477_ _3477_/A vssd1 vssd1 vccd1 vccd1 _6316_/D sky130_fd_sc_hd__clkbuf_1
X_5216_ _6311_/Q _6310_/Q _6309_/Q _6308_/Q vssd1 vssd1 vccd1 vccd1 _5218_/B sky130_fd_sc_hd__or4_1
XFILLER_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6196_ _6243_/A _6205_/B vssd1 vssd1 vccd1 vccd1 _6196_/X sky130_fd_sc_hd__or2_1
XFILLER_96_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5147_ _5160_/A _5147_/B _5147_/C vssd1 vssd1 vccd1 vccd1 _5148_/A sky130_fd_sc_hd__and3_1
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5078_ _6809_/Q _5078_/B vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__or2_1
X_4029_ _3986_/X _4028_/X _3633_/X vssd1 vssd1 vccd1 vccd1 _4029_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6869__129 vssd1 vssd1 vccd1 vccd1 _6869__129/HI _6978_/A sky130_fd_sc_hd__conb_1
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3400_ _6295_/Q _3396_/X _3398_/B vssd1 vssd1 vccd1 vccd1 _3400_/Y sky130_fd_sc_hd__a21boi_1
X_4380_ _4381_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3331_ _3331_/A _3331_/B _3331_/C _3331_/D vssd1 vssd1 vccd1 vccd1 _3332_/B sky130_fd_sc_hd__or4_4
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6050_ _6029_/X _6048_/X _6049_/X vssd1 vssd1 vccd1 vccd1 _6050_/X sky130_fd_sc_hd__a21o_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3262_/A vssd1 vssd1 vccd1 vccd1 _3262_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3193_ _3193_/A vssd1 vssd1 vccd1 vccd1 _3193_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5001_ _5001_/A vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__buf_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6952_ _6952_/A _3251_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
X_5903_ _5871_/X _5901_/X _5902_/X _5767_/X vssd1 vssd1 vccd1 vccd1 _5903_/X sky130_fd_sc_hd__a211o_1
X_5834_ _6713_/Q _5611_/X _5841_/S vssd1 vssd1 vccd1 vccd1 _5834_/X sky130_fd_sc_hd__mux2_1
X_5765_ _5765_/A _5765_/B vssd1 vssd1 vccd1 vccd1 _5765_/X sky130_fd_sc_hd__or2_1
X_4716_ _6371_/Q _4722_/B vssd1 vssd1 vccd1 vccd1 _4717_/A sky130_fd_sc_hd__and2_1
X_5696_ _6479_/Q _5678_/X _5680_/X _5693_/X _5695_/X vssd1 vssd1 vccd1 vccd1 _5696_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4647_ _4647_/A _4647_/B vssd1 vssd1 vccd1 vccd1 _6396_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4578_ _4597_/A _4595_/D _4579_/C vssd1 vssd1 vccd1 vccd1 _4580_/A sky130_fd_sc_hd__a21oi_1
X_6317_ _6523_/CLK _6317_/D vssd1 vssd1 vccd1 vccd1 _6317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3529_ _6651_/Q vssd1 vssd1 vccd1 vccd1 _3727_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6248_ _6248_/A vssd1 vssd1 vccd1 vccd1 _6248_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6179_ _6781_/Q _6169_/X _6177_/X _6178_/X vssd1 vssd1 vccd1 vccd1 _6781_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3880_ _3880_/A vssd1 vssd1 vccd1 vccd1 _6356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5550_ _6674_/Q _5523_/X _5547_/X _5549_/X _5540_/X vssd1 vssd1 vccd1 vccd1 _6674_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5481_ _5490_/A _5481_/B vssd1 vssd1 vccd1 vccd1 _5482_/A sky130_fd_sc_hd__and2_1
X_4501_ _4502_/B _4502_/C _4502_/A vssd1 vssd1 vccd1 vccd1 _4501_/Y sky130_fd_sc_hd__a21oi_2
X_4432_ _4576_/A _6374_/Q _6375_/Q _4510_/B vssd1 vssd1 vccd1 vccd1 _4436_/B sky130_fd_sc_hd__a22o_1
XANTENNA_0 _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4363_ _4363_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__xnor2_1
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3314_ _6494_/Q _6554_/Q vssd1 vssd1 vccd1 vccd1 _3370_/B sky130_fd_sc_hd__nor2b_2
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4294_ _6376_/Q vssd1 vssd1 vccd1 vccd1 _4393_/C sky130_fd_sc_hd__clkbuf_2
X_6102_ _6102_/A vssd1 vssd1 vccd1 vccd1 _6102_/X sky130_fd_sc_hd__clkbuf_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3249_/A vssd1 vssd1 vccd1 vccd1 _3245_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6033_ _6029_/X _6030_/X _6032_/X vssd1 vssd1 vccd1 vccd1 _6033_/X sky130_fd_sc_hd__a21o_1
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6935_ _6935_/A _3230_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6797_ _6799_/CLK _6797_/D vssd1 vssd1 vccd1 vccd1 _6797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5817_ _6709_/Q _5797_/X _5816_/X _5810_/X vssd1 vssd1 vccd1 vccd1 _6709_/D sky130_fd_sc_hd__o211a_1
X_5748_ _5619_/X _5698_/X _5699_/X _5747_/X vssd1 vssd1 vccd1 vccd1 _5748_/X sky130_fd_sc_hd__o211a_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5679_ _5957_/C _6062_/C vssd1 vssd1 vccd1 vccd1 _5735_/A sky130_fd_sc_hd__nand2_2
XFILLER_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _6544_/Q _4982_/B vssd1 vssd1 vccd1 vccd1 _4986_/B sky130_fd_sc_hd__and2_1
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6720_ _6799_/CLK _6720_/D vssd1 vssd1 vccd1 vccd1 _6720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3932_ _3933_/A _3933_/B vssd1 vssd1 vccd1 vccd1 _3934_/B sky130_fd_sc_hd__nand2_1
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6651_ _6763_/CLK _6651_/D vssd1 vssd1 vccd1 vccd1 _6651_/Q sky130_fd_sc_hd__dfxtp_1
X_3863_ _3860_/A _3862_/X _3340_/X vssd1 vssd1 vccd1 vccd1 _6349_/D sky130_fd_sc_hd__o21a_1
X_6582_ _6586_/CLK _6582_/D vssd1 vssd1 vccd1 vccd1 _6920_/A sky130_fd_sc_hd__dfxtp_1
X_5602_ _6470_/Q vssd1 vssd1 vccd1 vccd1 _5602_/X sky130_fd_sc_hd__buf_2
XFILLER_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3794_ _3764_/A _3763_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3795_/B sky130_fd_sc_hd__o21ba_1
X_5533_ _6479_/Q vssd1 vssd1 vccd1 vccd1 _6233_/A sky130_fd_sc_hd__buf_4
X_5464_ _5474_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _5465_/A sky130_fd_sc_hd__and2_1
X_5395_ _5395_/A vssd1 vssd1 vccd1 vccd1 _6639_/D sky130_fd_sc_hd__clkbuf_1
X_4415_ _4414_/B _4414_/C _4414_/A vssd1 vssd1 vccd1 vccd1 _4416_/C sky130_fd_sc_hd__o21ai_1
XFILLER_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4346_ _4381_/A vssd1 vssd1 vccd1 vccd1 _4348_/A sky130_fd_sc_hd__inv_2
XFILLER_113_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4277_ _6664_/Q vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3228_ _3231_/A vssd1 vssd1 vccd1 vccd1 _3228_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6016_ _6743_/Q _6011_/X _6015_/X _5999_/X vssd1 vssd1 vccd1 vccd1 _6743_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _6918_/A _3210_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__ebufn_8
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ _4227_/A _4228_/A _4270_/A _4230_/C vssd1 vssd1 vccd1 vccd1 _4201_/B sky130_fd_sc_hd__nand4_1
X_5180_ _6919_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5184_/B sky130_fd_sc_hd__or2_1
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4131_ _4144_/B _4144_/C _4144_/A vssd1 vssd1 vccd1 vccd1 _4131_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4062_ _4062_/A _4062_/B _4062_/C vssd1 vssd1 vccd1 vccd1 _4062_/X sky130_fd_sc_hd__and3_2
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4964_ _4969_/C _5239_/B _4964_/C vssd1 vssd1 vccd1 vccd1 _4965_/A sky130_fd_sc_hd__and3b_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6703_ _6809_/CLK _6703_/D vssd1 vssd1 vccd1 vccd1 _6703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3915_ _3915_/A vssd1 vssd1 vccd1 vccd1 _6360_/D sky130_fd_sc_hd__clkbuf_1
X_4895_ _4895_/A vssd1 vssd1 vccd1 vccd1 _4895_/X sky130_fd_sc_hd__clkbuf_2
X_6634_ _6532_/Q _6634_/D vssd1 vssd1 vccd1 vccd1 _6634_/Q sky130_fd_sc_hd__dfxtp_1
X_3846_ _3827_/X _3828_/X _3843_/Y _3825_/Y vssd1 vssd1 vccd1 vccd1 _3846_/X sky130_fd_sc_hd__a211o_1
XFILLER_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6565_ _6569_/CLK _6565_/D vssd1 vssd1 vccd1 vccd1 _6903_/A sky130_fd_sc_hd__dfxtp_1
X_3777_ _3826_/B _3777_/B vssd1 vssd1 vccd1 vccd1 _3828_/B sky130_fd_sc_hd__or2_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6496_ _6528_/CLK _6496_/D hold3/X vssd1 vssd1 vccd1 vccd1 _6496_/Q sky130_fd_sc_hd__dfrtp_1
X_5516_ _5922_/A vssd1 vssd1 vccd1 vccd1 _5638_/A sky130_fd_sc_hd__clkbuf_4
X_5447_ _5447_/A vssd1 vssd1 vccd1 vccd1 _6656_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5378_ _5378_/A vssd1 vssd1 vccd1 vccd1 _6635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4329_ _6378_/Q vssd1 vssd1 vccd1 vccd1 _4576_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _3596_/A _3810_/B _3653_/B _3698_/Y vssd1 vssd1 vccd1 vccd1 _3701_/B sky130_fd_sc_hd__a211oi_1
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4680_ _6347_/Q _4688_/B vssd1 vssd1 vccd1 vccd1 _4681_/A sky130_fd_sc_hd__and2_1
XFILLER_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3631_ _3629_/X _3631_/B vssd1 vssd1 vccd1 vccd1 _3631_/X sky130_fd_sc_hd__and2b_1
X_3562_ _3563_/A _3563_/B vssd1 vssd1 vccd1 vccd1 _3568_/A sky130_fd_sc_hd__or2_1
X_6350_ _6763_/CLK _6350_/D vssd1 vssd1 vccd1 vccd1 _6350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5301_ _6614_/Q _5305_/B vssd1 vssd1 vccd1 vccd1 _5302_/A sky130_fd_sc_hd__and2_1
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3493_ _6324_/Q _6528_/Q _3495_/S vssd1 vssd1 vccd1 vccd1 _3494_/A sky130_fd_sc_hd__mux2_1
X_6281_ _6268_/X _6280_/Y _6264_/X vssd1 vssd1 vccd1 vccd1 _6281_/Y sky130_fd_sc_hd__o21ai_1
X_5232_ _6608_/Q _6607_/Q _5232_/C vssd1 vssd1 vccd1 vccd1 _5414_/C sky130_fd_sc_hd__or3_1
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5163_ _6916_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5166_/B sky130_fd_sc_hd__or2_1
XFILLER_110_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4114_ _4153_/A _4153_/B _4114_/C _4153_/C vssd1 vssd1 vccd1 vccd1 _4156_/A sky130_fd_sc_hd__nand4_2
XFILLER_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5094_ _5081_/X _5092_/X _5093_/X _5088_/X vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__a31o_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4045_ _4083_/A _4151_/B vssd1 vssd1 vccd1 vccd1 _4093_/A sky130_fd_sc_hd__nand2_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _6023_/A vssd1 vssd1 vccd1 vccd1 _5996_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4947_ _4950_/B _4945_/X _4946_/Y vssd1 vssd1 vccd1 vccd1 _6533_/D sky130_fd_sc_hd__o21a_1
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4878_ _6504_/Q _4870_/X _4873_/X input62/X vssd1 vssd1 vccd1 vccd1 _6504_/D sky130_fd_sc_hd__a22o_1
X_6617_ _6667_/CLK _6617_/D vssd1 vssd1 vccd1 vccd1 _6617_/Q sky130_fd_sc_hd__dfxtp_1
X_3829_ _3825_/Y _3827_/X _3828_/X _3636_/A vssd1 vssd1 vccd1 vccd1 _3829_/X sky130_fd_sc_hd__a31o_1
XFILLER_116_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6548_ _6551_/CLK _6548_/D vssd1 vssd1 vccd1 vccd1 _6548_/Q sky130_fd_sc_hd__dfxtp_1
X_6479_ _6763_/CLK _6479_/D vssd1 vssd1 vccd1 vccd1 _6479_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6817__77 vssd1 vssd1 vccd1 vccd1 _6817__77/HI _6926_/A sky130_fd_sc_hd__conb_1
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6831__91 vssd1 vssd1 vccd1 vccd1 _6831__91/HI _6940_/A sky130_fd_sc_hd__conb_1
XFILLER_0_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5850_ _5946_/A vssd1 vssd1 vccd1 vccd1 _5850_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5781_ _6632_/Q _6631_/Q _5971_/A _6629_/Q vssd1 vssd1 vccd1 vccd1 _5872_/B sky130_fd_sc_hd__or4b_1
X_4801_ _4801_/A vssd1 vssd1 vccd1 vccd1 _6465_/D sky130_fd_sc_hd__clkbuf_1
X_4732_ _4732_/A vssd1 vssd1 vccd1 vccd1 _6434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4663_ _4663_/A vssd1 vssd1 vccd1 vccd1 _6403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3614_ _3614_/A _3614_/B _3614_/C vssd1 vssd1 vccd1 vccd1 _3622_/B sky130_fd_sc_hd__nand3_2
X_6402_ _6789_/CLK _6402_/D vssd1 vssd1 vccd1 vccd1 _6402_/Q sky130_fd_sc_hd__dfxtp_1
X_4594_ _4622_/A _4595_/C _4595_/D _4623_/A vssd1 vssd1 vccd1 vccd1 _4596_/A sky130_fd_sc_hd__a22o_1
X_6333_ _6551_/CLK _6333_/D vssd1 vssd1 vccd1 vccd1 _6333_/Q sky130_fd_sc_hd__dfxtp_1
X_3545_ _3899_/A _3545_/B _3565_/B vssd1 vssd1 vccd1 vccd1 _3546_/A sky130_fd_sc_hd__and3_1
XFILLER_115_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6264_ _6264_/A vssd1 vssd1 vccd1 vccd1 _6264_/X sky130_fd_sc_hd__buf_2
X_3476_ _6316_/Q _6520_/Q _3484_/S vssd1 vssd1 vccd1 vccd1 _3477_/A sky130_fd_sc_hd__mux2_1
X_5215_ _6307_/Q _6306_/Q _6305_/Q _6304_/Q vssd1 vssd1 vccd1 vccd1 _5218_/A sky130_fd_sc_hd__or4_1
X_6195_ _6222_/B vssd1 vssd1 vccd1 vccd1 _6205_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5146_ _5119_/X _5144_/X _5145_/X vssd1 vssd1 vccd1 vccd1 _5147_/C sky130_fd_sc_hd__a21o_1
XFILLER_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5077_ _5077_/A _5077_/B vssd1 vssd1 vccd1 vccd1 _5077_/X sky130_fd_sc_hd__or2_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4028_ _4026_/X _4028_/B vssd1 vssd1 vccd1 vccd1 _4028_/X sky130_fd_sc_hd__and2b_1
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5979_ _6736_/Q _5946_/X _5978_/X _5959_/X vssd1 vssd1 vccd1 vccd1 _6736_/D sky130_fd_sc_hd__o211a_1
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3330_ _3330_/A _3330_/B _3330_/C _3330_/D vssd1 vssd1 vccd1 vccd1 _3332_/A sky130_fd_sc_hd__or4_1
XFILLER_112_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5000_ _5000_/A vssd1 vssd1 vccd1 vccd1 _6549_/D sky130_fd_sc_hd__clkbuf_1
X_3261_ _3262_/A vssd1 vssd1 vccd1 vccd1 _3261_/Y sky130_fd_sc_hd__inv_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3192_ _3193_/A vssd1 vssd1 vccd1 vccd1 _3192_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6951_ _6951_/A _3249_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5902_ _6482_/Q _5964_/D _5914_/C vssd1 vssd1 vccd1 vccd1 _5902_/X sky130_fd_sc_hd__and3_1
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5833_ _6712_/Q _5825_/X _5832_/X _5810_/X vssd1 vssd1 vccd1 vccd1 _6712_/D sky130_fd_sc_hd__o211a_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6852__112 vssd1 vssd1 vccd1 vccd1 _6852__112/HI _6961_/A sky130_fd_sc_hd__conb_1
X_5764_ _6702_/Q _5660_/X _5764_/S vssd1 vssd1 vccd1 vccd1 _5765_/B sky130_fd_sc_hd__mux2_1
X_4715_ _4715_/A vssd1 vssd1 vccd1 vccd1 _6426_/D sky130_fd_sc_hd__clkbuf_1
X_5695_ _5915_/A vssd1 vssd1 vccd1 vccd1 _5695_/X sky130_fd_sc_hd__clkbuf_2
X_4646_ _4644_/X _4633_/X _4635_/Y _4385_/A vssd1 vssd1 vccd1 vccd1 _4647_/B sky130_fd_sc_hd__a31o_1
X_4577_ _4577_/A _4600_/A vssd1 vssd1 vccd1 vccd1 _4579_/C sky130_fd_sc_hd__nor2_1
X_6316_ _6523_/CLK _6316_/D vssd1 vssd1 vccd1 vccd1 _6316_/Q sky130_fd_sc_hd__dfxtp_1
X_3528_ _3528_/A vssd1 vssd1 vccd1 vccd1 _6336_/D sky130_fd_sc_hd__clkbuf_1
X_3459_ _3459_/A vssd1 vssd1 vccd1 vccd1 _6308_/D sky130_fd_sc_hd__clkbuf_1
X_6247_ _6267_/A vssd1 vssd1 vccd1 vccd1 _6247_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6178_ _6178_/A vssd1 vssd1 vccd1 vccd1 _6178_/X sky130_fd_sc_hd__buf_2
XFILLER_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5129_ _5129_/A _5129_/B _5129_/C vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__and3_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5480_ _6314_/Q _4333_/A _5483_/S vssd1 vssd1 vccd1 vccd1 _5481_/B sky130_fd_sc_hd__mux2_1
X_4500_ _4283_/A _4637_/B _4453_/B _4499_/X vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__a31o_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_1 _5081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4431_ _6670_/Q vssd1 vssd1 vccd1 vccd1 _4510_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4362_ _4449_/A _4595_/C vssd1 vssd1 vccd1 vccd1 _4363_/B sky130_fd_sc_hd__nand2_1
X_4293_ _4293_/A vssd1 vssd1 vccd1 vccd1 _6383_/D sky130_fd_sc_hd__clkbuf_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3313_/Y sky130_fd_sc_hd__inv_2
X_6101_ _6469_/Q _6081_/X _6096_/X _6087_/X _6485_/Q vssd1 vssd1 vccd1 vccd1 _6101_/X
+ sky130_fd_sc_hd__a32o_1
X_3244_ _3250_/A vssd1 vssd1 vccd1 vccd1 _3249_/A sky130_fd_sc_hd__buf_8
XFILLER_112_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6032_ _6488_/Q _6023_/X _6013_/X _6031_/X vssd1 vssd1 vccd1 vccd1 _6032_/X sky130_fd_sc_hd__a31o_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6934_ _6934_/A _3229_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6796_ _6799_/CLK _6796_/D vssd1 vssd1 vccd1 vccd1 _6796_/Q sky130_fd_sc_hd__dfxtp_1
X_5816_ _6483_/Q _5812_/X _5814_/X _5808_/X _5815_/X vssd1 vssd1 vccd1 vccd1 _5816_/X
+ sky130_fd_sc_hd__a221o_1
X_5747_ _5765_/A _5747_/B vssd1 vssd1 vccd1 vccd1 _5747_/X sky130_fd_sc_hd__or2_1
XFILLER_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5678_ _5734_/A vssd1 vssd1 vccd1 vccd1 _5678_/X sky130_fd_sc_hd__clkbuf_2
X_4629_ _4642_/B _4629_/B vssd1 vssd1 vccd1 vccd1 _4630_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4980_ _6333_/Q _4980_/B _4993_/A _5008_/C vssd1 vssd1 vccd1 vccd1 _4982_/B sky130_fd_sc_hd__and4_1
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3931_ _3953_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _3933_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6650_ _6763_/CLK _6650_/D vssd1 vssd1 vccd1 vccd1 _6650_/Q sky130_fd_sc_hd__dfxtp_1
X_3862_ _3850_/A _3881_/A _3861_/X _3857_/A vssd1 vssd1 vccd1 vccd1 _3862_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6581_ _6586_/CLK _6581_/D vssd1 vssd1 vccd1 vccd1 _6919_/A sky130_fd_sc_hd__dfxtp_1
X_5601_ _5650_/A vssd1 vssd1 vccd1 vccd1 _5601_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3793_ _3793_/A _3813_/B vssd1 vssd1 vccd1 vccd1 _3815_/B sky130_fd_sc_hd__nor2_1
X_5532_ _5524_/X _5525_/X _5505_/X _5531_/X vssd1 vssd1 vccd1 vccd1 _5532_/X sky130_fd_sc_hd__o211a_1
X_5463_ _6309_/Q _4202_/A _5466_/S vssd1 vssd1 vccd1 vccd1 _5464_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5394_ _6639_/Q _5396_/B vssd1 vssd1 vccd1 vccd1 _5395_/A sky130_fd_sc_hd__and2_1
X_4414_ _4414_/A _4414_/B _4414_/C vssd1 vssd1 vccd1 vccd1 _4416_/B sky130_fd_sc_hd__or3_2
XFILLER_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4345_ _4347_/A _4347_/B vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4276_ _4276_/A vssd1 vssd1 vccd1 vccd1 _6381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6015_ _6001_/X _6012_/X _6014_/X vssd1 vssd1 vccd1 vccd1 _6015_/X sky130_fd_sc_hd__a21o_1
X_3227_ _3231_/A vssd1 vssd1 vccd1 vccd1 _3227_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6917_ _6917_/A _3209_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__ebufn_8
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6779_ _6532_/Q _6779_/D vssd1 vssd1 vccd1 vccd1 _6779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4130_ _3941_/A _4230_/C _4087_/B _4086_/B vssd1 vssd1 vccd1 vccd1 _4144_/A sky130_fd_sc_hd__a31o_1
XFILLER_122_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4061_ _4062_/B _4062_/C _4062_/A vssd1 vssd1 vccd1 vccd1 _4061_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4963_ _4962_/B _4962_/C _6538_/Q vssd1 vssd1 vccd1 vccd1 _4964_/C sky130_fd_sc_hd__a21o_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6702_ _6809_/CLK _6702_/D vssd1 vssd1 vccd1 vccd1 _6702_/Q sky130_fd_sc_hd__dfxtp_1
X_3914_ _4325_/A _3914_/B _3933_/A vssd1 vssd1 vccd1 vccd1 _3915_/A sky130_fd_sc_hd__and3_1
X_4894_ _4910_/S vssd1 vssd1 vccd1 vccd1 _4894_/X sky130_fd_sc_hd__clkbuf_2
X_6633_ _6532_/Q _6633_/D vssd1 vssd1 vccd1 vccd1 _6633_/Q sky130_fd_sc_hd__dfxtp_1
X_3845_ _3847_/A _3831_/B _3843_/Y _3844_/Y _3633_/X vssd1 vssd1 vccd1 vccd1 _6347_/D
+ sky130_fd_sc_hd__a311oi_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6564_ _6569_/CLK _6564_/D vssd1 vssd1 vccd1 vccd1 _6902_/A sky130_fd_sc_hd__dfxtp_1
X_3776_ _3826_/A _3775_/B _3775_/C vssd1 vssd1 vccd1 vccd1 _3777_/B sky130_fd_sc_hd__o21a_1
X_6495_ _6554_/CLK _6495_/D hold3/A vssd1 vssd1 vccd1 vccd1 _6495_/Q sky130_fd_sc_hd__dfrtp_2
X_5515_ _5506_/X _5512_/X _5631_/A vssd1 vssd1 vccd1 vccd1 _5515_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5446_ _5456_/A _5446_/B vssd1 vssd1 vccd1 vccd1 _5447_/A sky130_fd_sc_hd__and2_1
X_5377_ _6635_/Q _5396_/B vssd1 vssd1 vccd1 vccd1 _5378_/A sky130_fd_sc_hd__and2_1
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4328_ _4354_/C _4328_/B vssd1 vssd1 vccd1 vccd1 _4332_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4259_ _4259_/A vssd1 vssd1 vccd1 vccd1 _5458_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3630_ _3629_/A _3629_/B _3629_/C vssd1 vssd1 vccd1 vccd1 _3631_/B sky130_fd_sc_hd__a21o_1
X_3561_ _3534_/Y _3549_/B _3538_/B _3538_/A vssd1 vssd1 vccd1 vccd1 _3563_/B sky130_fd_sc_hd__o22a_1
X_5300_ _5300_/A vssd1 vssd1 vccd1 vccd1 _6613_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3492_ _3492_/A vssd1 vssd1 vccd1 vccd1 _6323_/D sky130_fd_sc_hd__clkbuf_1
X_6280_ _6280_/A _6283_/B vssd1 vssd1 vccd1 vccd1 _6280_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5231_ _6600_/Q _6599_/Q _6595_/Q _6592_/Q vssd1 vssd1 vccd1 vccd1 _5232_/C sky130_fd_sc_hd__or4_1
XFILLER_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5162_ _5162_/A vssd1 vssd1 vccd1 vccd1 _5191_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5093_ _6811_/Q _5109_/B vssd1 vssd1 vccd1 vccd1 _5093_/X sky130_fd_sc_hd__or2_1
X_4113_ _6663_/Q _6352_/Q _6353_/Q _4153_/B vssd1 vssd1 vccd1 vccd1 _4116_/C sky130_fd_sc_hd__a22o_1
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4044_ _4043_/B _4043_/C _4043_/A vssd1 vssd1 vccd1 vccd1 _4052_/C sky130_fd_sc_hd__a21o_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5995_ _6740_/Q _5560_/X _6017_/S vssd1 vssd1 vccd1 vccd1 _5995_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4946_ _4950_/B _5041_/A _3637_/A vssd1 vssd1 vccd1 vccd1 _4946_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4877_ _6503_/Q _4870_/X _4873_/X input61/X vssd1 vssd1 vccd1 vccd1 _6503_/D sky130_fd_sc_hd__a22o_1
X_6616_ _6667_/CLK _6616_/D vssd1 vssd1 vccd1 vccd1 _6616_/Q sky130_fd_sc_hd__dfxtp_1
X_3828_ _3828_/A _3828_/B _3828_/C _3828_/D vssd1 vssd1 vccd1 vccd1 _3828_/X sky130_fd_sc_hd__or4_2
X_6547_ _6551_/CLK _6547_/D vssd1 vssd1 vccd1 vccd1 _6547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3759_ _3759_/A vssd1 vssd1 vccd1 vccd1 _3835_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6478_ _6795_/CLK _6478_/D vssd1 vssd1 vccd1 vccd1 _6478_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5429_ _5439_/A _5429_/B vssd1 vssd1 vccd1 vccd1 _5430_/A sky130_fd_sc_hd__and2_1
XFILLER_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6522_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4800_ _6417_/Q _4800_/B vssd1 vssd1 vccd1 vccd1 _4801_/A sky130_fd_sc_hd__and2_1
XFILLER_22_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5780_ _6704_/Q _5508_/X _5859_/S vssd1 vssd1 vccd1 vccd1 _5780_/X sky130_fd_sc_hd__mux2_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _6386_/Q _4733_/B vssd1 vssd1 vccd1 vccd1 _4732_/A sky130_fd_sc_hd__and2_1
X_4662_ _6339_/Q _4666_/B vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__and2_1
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3613_ _3641_/A _3660_/B _3641_/C vssd1 vssd1 vccd1 vccd1 _3614_/C sky130_fd_sc_hd__a21o_1
X_6401_ _6789_/CLK _6401_/D vssd1 vssd1 vccd1 vccd1 _6401_/Q sky130_fd_sc_hd__dfxtp_1
X_4593_ _4593_/A _4593_/B vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__or2_1
X_6332_ _6551_/CLK _6332_/D vssd1 vssd1 vccd1 vccd1 _6332_/Q sky130_fd_sc_hd__dfxtp_1
X_3544_ _3544_/A _3544_/B vssd1 vssd1 vccd1 vccd1 _3565_/B sky130_fd_sc_hd__or2_1
X_3475_ _3486_/A vssd1 vssd1 vccd1 vccd1 _3484_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6263_ _6263_/A _6263_/B vssd1 vssd1 vccd1 vccd1 _6263_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5214_ _5214_/A _5214_/B _5214_/C _5214_/D vssd1 vssd1 vccd1 vccd1 _5224_/A sky130_fd_sc_hd__or4_4
X_6194_ _6207_/A vssd1 vssd1 vccd1 vccd1 _6194_/X sky130_fd_sc_hd__buf_2
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5145_ _5176_/A vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _6681_/Q _6713_/Q _6745_/Q _6777_/Q _5049_/X _5063_/X vssd1 vssd1 vccd1 vccd1
+ _5077_/B sky130_fd_sc_hd__mux4_1
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4027_ _4026_/A _4026_/B _4026_/C vssd1 vssd1 vccd1 vccd1 _4028_/B sky130_fd_sc_hd__a21o_1
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _5969_/X _5974_/X _5977_/X vssd1 vssd1 vccd1 vccd1 _5978_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ _4928_/X _6531_/Q _4929_/S vssd1 vssd1 vccd1 vccd1 _4930_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3262_/A vssd1 vssd1 vccd1 vccd1 _3260_/Y sky130_fd_sc_hd__inv_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3193_/A vssd1 vssd1 vccd1 vccd1 _3191_/Y sky130_fd_sc_hd__inv_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6950_ _6950_/A _3248_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5901_ _5560_/X _5889_/X _5891_/X _5874_/X _6724_/Q vssd1 vssd1 vccd1 vccd1 _5901_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5832_ _6486_/Q _5812_/X _5831_/X _5808_/X _5815_/X vssd1 vssd1 vccd1 vccd1 _5832_/X
+ sky130_fd_sc_hd__a221o_1
X_6891__151 vssd1 vssd1 vccd1 vccd1 _6891__151/HI _7000_/A sky130_fd_sc_hd__conb_1
X_5763_ _6701_/Q _5755_/X _5762_/X _5739_/X vssd1 vssd1 vccd1 vccd1 _6701_/D sky130_fd_sc_hd__o211a_1
X_4714_ _6370_/Q _4722_/B vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__and2_1
X_5694_ _6031_/A vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__clkbuf_2
X_4645_ _4633_/X _4635_/Y _4644_/X vssd1 vssd1 vccd1 vccd1 _4647_/A sky130_fd_sc_hd__a21oi_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4576_ _4576_/A _4576_/B _4576_/C _6379_/Q vssd1 vssd1 vccd1 vccd1 _4600_/A sky130_fd_sc_hd__and4_1
X_6315_ _6531_/CLK _6315_/D vssd1 vssd1 vccd1 vccd1 _6315_/Q sky130_fd_sc_hd__dfxtp_1
X_3527_ _3899_/A _3527_/B _3544_/A vssd1 vssd1 vccd1 vccd1 _3528_/A sky130_fd_sc_hd__and3_1
XFILLER_103_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3458_ _6308_/Q _6512_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _3459_/A sky130_fd_sc_hd__mux2_1
X_6246_ _6804_/Q _6226_/X _6245_/Y _6235_/X vssd1 vssd1 vccd1 vccd1 _6804_/D sky130_fd_sc_hd__o211a_1
X_3389_ _6291_/Q _3390_/C _3388_/Y vssd1 vssd1 vccd1 vccd1 _6291_/D sky130_fd_sc_hd__a21oi_1
X_6177_ _6280_/A _6180_/B vssd1 vssd1 vccd1 vccd1 _6177_/X sky130_fd_sc_hd__or2_1
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5128_ _5119_/X _5127_/X _5115_/X vssd1 vssd1 vccd1 vccd1 _5129_/C sky130_fd_sc_hd__a21o_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5059_ _5077_/A _5059_/B vssd1 vssd1 vccd1 vccd1 _5059_/X sky130_fd_sc_hd__or2_1
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6875__135 vssd1 vssd1 vccd1 vccd1 _6875__135/HI _6984_/A sky130_fd_sc_hd__conb_1
XFILLER_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4430_ _6671_/Q vssd1 vssd1 vccd1 vccd1 _4576_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_2 _5552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _4547_/B vssd1 vssd1 vccd1 vccd1 _4595_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6100_ _6100_/A vssd1 vssd1 vccd1 vccd1 _6758_/D sky130_fd_sc_hd__clkbuf_1
X_3312_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3312_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4292_ _4325_/A _4292_/B _4304_/A vssd1 vssd1 vccd1 vccd1 _4293_/A sky130_fd_sc_hd__and3_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _6031_/A vssd1 vssd1 vccd1 vccd1 _6031_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3243_/A vssd1 vssd1 vccd1 vccd1 _3243_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6933_ _6933_/A _3228_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_81_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5815_ _5843_/A vssd1 vssd1 vccd1 vccd1 _5815_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6795_ _6795_/CLK _6795_/D vssd1 vssd1 vccd1 vccd1 _6795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5746_ _6698_/Q _5621_/X _5764_/S vssd1 vssd1 vccd1 vccd1 _5747_/B sky130_fd_sc_hd__mux2_1
X_5677_ _5870_/B _6062_/C vssd1 vssd1 vccd1 vccd1 _5734_/A sky130_fd_sc_hd__and2b_2
X_4628_ _4638_/A _4642_/A vssd1 vssd1 vccd1 vccd1 _4629_/B sky130_fd_sc_hd__nor2_1
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4559_ _4572_/A _4557_/X _4518_/B _4541_/Y vssd1 vssd1 vccd1 vccd1 _4559_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6229_ _6229_/A _6243_/B vssd1 vssd1 vccd1 vccd1 _6229_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6859__119 vssd1 vssd1 vccd1 vccd1 _6859__119/HI _6968_/A sky130_fd_sc_hd__conb_1
XFILLER_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3930_ _3930_/A _3930_/B vssd1 vssd1 vccd1 vccd1 _3931_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _3849_/A _3879_/A _3853_/B vssd1 vssd1 vccd1 vccd1 _3861_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6580_ _6580_/CLK _6580_/D vssd1 vssd1 vccd1 vccd1 _6918_/A sky130_fd_sc_hd__dfxtp_1
X_3792_ _3810_/A _3792_/B _3792_/C vssd1 vssd1 vccd1 vccd1 _3813_/B sky130_fd_sc_hd__and3_1
X_5600_ _6679_/Q _5551_/X _5597_/X _5599_/X _5591_/X vssd1 vssd1 vccd1 vccd1 _6679_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5531_ _5575_/A _5531_/B vssd1 vssd1 vccd1 vccd1 _5531_/X sky130_fd_sc_hd__or2_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5462_ _5462_/A vssd1 vssd1 vccd1 vccd1 _6660_/D sky130_fd_sc_hd__clkbuf_1
X_4413_ _4428_/A _4428_/B _4428_/C vssd1 vssd1 vccd1 vccd1 _4414_/C sky130_fd_sc_hd__and3_1
X_5393_ _5393_/A vssd1 vssd1 vccd1 vccd1 _6638_/D sky130_fd_sc_hd__clkbuf_1
X_4344_ _4354_/B _4315_/X _4320_/A vssd1 vssd1 vccd1 vccd1 _4347_/B sky130_fd_sc_hd__a21o_1
XFILLER_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4275_ _4275_/A _4655_/B vssd1 vssd1 vccd1 vccd1 _4276_/A sky130_fd_sc_hd__and2_1
X_6014_ _6485_/Q _5996_/X _6013_/X _6003_/X vssd1 vssd1 vccd1 vccd1 _6014_/X sky130_fd_sc_hd__a31o_1
X_3226_ _3250_/A vssd1 vssd1 vccd1 vccd1 _3231_/A sky130_fd_sc_hd__buf_12
XFILLER_55_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6916_ _6916_/A _3208_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__ebufn_8
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6546_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_6778_ _6532_/Q _6778_/D vssd1 vssd1 vccd1 vccd1 _6778_/Q sky130_fd_sc_hd__dfxtp_1
X_5729_ _6695_/Q _5594_/X _5751_/S vssd1 vssd1 vccd1 vccd1 _5729_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6838__98 vssd1 vssd1 vccd1 vccd1 _6838__98/HI _6947_/A sky130_fd_sc_hd__conb_1
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4060_ _4060_/A _4060_/B vssd1 vssd1 vccd1 vccd1 _4062_/A sky130_fd_sc_hd__xnor2_1
XFILLER_37_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4962_ _6538_/Q _4962_/B _4962_/C vssd1 vssd1 vccd1 vccd1 _4969_/C sky130_fd_sc_hd__and3_1
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6701_ _6799_/CLK _6701_/D vssd1 vssd1 vccd1 vccd1 _6701_/Q sky130_fd_sc_hd__dfxtp_1
X_4893_ _6514_/Q _4887_/X _4888_/X input41/X vssd1 vssd1 vccd1 vccd1 _6514_/D sky130_fd_sc_hd__a22o_1
X_3913_ _3913_/A _3928_/B _3911_/X vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__or3b_1
X_6632_ _6799_/CLK _6632_/D vssd1 vssd1 vccd1 vccd1 _6632_/Q sky130_fd_sc_hd__dfxtp_1
X_3844_ _3847_/A _3831_/B _3843_/Y vssd1 vssd1 vccd1 vccd1 _3844_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6563_ _6569_/CLK _6563_/D vssd1 vssd1 vccd1 vccd1 _6901_/A sky130_fd_sc_hd__dfxtp_1
X_3775_ _3826_/A _3775_/B _3775_/C vssd1 vssd1 vccd1 vccd1 _3826_/B sky130_fd_sc_hd__nor3_1
XFILLER_20_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6494_ _6554_/CLK _6494_/D hold3/A vssd1 vssd1 vccd1 vccd1 _6494_/Q sky130_fd_sc_hd__dfrtp_1
X_5514_ _5873_/A _5700_/A vssd1 vssd1 vccd1 vccd1 _5631_/A sky130_fd_sc_hd__or2_2
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5445_ _6304_/Q _3889_/A _5448_/S vssd1 vssd1 vccd1 vccd1 _5446_/B sky130_fd_sc_hd__mux2_1
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5376_ _5376_/A vssd1 vssd1 vccd1 vccd1 _6634_/D sky130_fd_sc_hd__clkbuf_1
X_4327_ _6665_/Q _4354_/B vssd1 vssd1 vccd1 vccd1 _4328_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4258_ _4258_/A vssd1 vssd1 vccd1 vccd1 _6374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3209_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3209_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4189_ _4189_/A _4157_/A vssd1 vssd1 vccd1 vccd1 _4189_/X sky130_fd_sc_hd__or2b_1
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3560_ _3571_/A _3571_/B vssd1 vssd1 vccd1 vccd1 _3563_/A sky130_fd_sc_hd__xnor2_1
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5230_ _6611_/Q _6610_/Q _5230_/C _5230_/D vssd1 vssd1 vccd1 vccd1 _5236_/B sky130_fd_sc_hd__nor4_1
X_3491_ _6323_/Q _6527_/Q _3495_/S vssd1 vssd1 vccd1 vccd1 _3492_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5161_ _5161_/A vssd1 vssd1 vccd1 vccd1 _6577_/D sky130_fd_sc_hd__clkbuf_1
X_5092_ _5108_/A _5092_/B vssd1 vssd1 vccd1 vccd1 _5092_/X sky130_fd_sc_hd__or2_1
X_4112_ _4109_/X _4220_/A _4111_/Y vssd1 vssd1 vccd1 vccd1 _6366_/D sky130_fd_sc_hd__a21oi_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4043_ _4043_/A _4043_/B _4043_/C vssd1 vssd1 vccd1 vccd1 _4052_/B sky130_fd_sc_hd__nand3_1
XFILLER_77_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5994_ _6048_/S vssd1 vssd1 vccd1 vccd1 _6017_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4945_ _5041_/A vssd1 vssd1 vccd1 vccd1 _4945_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _6502_/Q _4870_/X _4873_/X input58/X vssd1 vssd1 vccd1 vccd1 _6502_/D sky130_fd_sc_hd__a22o_1
X_6615_ _6667_/CLK _6615_/D vssd1 vssd1 vccd1 vccd1 _6615_/Q sky130_fd_sc_hd__dfxtp_1
X_3827_ _3828_/B _3779_/X _3828_/D _3826_/Y _3803_/B vssd1 vssd1 vccd1 vccd1 _3827_/X
+ sky130_fd_sc_hd__o32a_1
X_6546_ _6546_/CLK _6546_/D vssd1 vssd1 vccd1 vccd1 _6546_/Q sky130_fd_sc_hd__dfxtp_1
X_3758_ _3810_/A _3758_/B vssd1 vssd1 vccd1 vccd1 _3764_/A sky130_fd_sc_hd__nand2_1
X_6477_ _6763_/CLK _6477_/D vssd1 vssd1 vccd1 vccd1 _6477_/Q sky130_fd_sc_hd__dfxtp_2
X_3689_ _3690_/B _3789_/C _3605_/B _3753_/A vssd1 vssd1 vccd1 vccd1 _3691_/A sky130_fd_sc_hd__a22oi_1
X_5428_ _5217_/A _3755_/B _5431_/S vssd1 vssd1 vccd1 vccd1 _5429_/B sky130_fd_sc_hd__mux2_1
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5359_ _5882_/A vssd1 vssd1 vccd1 vccd1 _5873_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4730_/A vssd1 vssd1 vccd1 vccd1 _6433_/D sky130_fd_sc_hd__clkbuf_1
X_4661_ _4661_/A vssd1 vssd1 vccd1 vccd1 _6402_/D sky130_fd_sc_hd__clkbuf_1
X_3612_ _3641_/A _3660_/B _3641_/C vssd1 vssd1 vccd1 vccd1 _3614_/B sky130_fd_sc_hd__nand3_1
X_6400_ _6789_/CLK _6400_/D vssd1 vssd1 vccd1 vccd1 _6400_/Q sky130_fd_sc_hd__dfxtp_1
X_6331_ _6546_/CLK _6331_/D vssd1 vssd1 vccd1 vccd1 _6331_/Q sky130_fd_sc_hd__dfxtp_1
X_4592_ _4990_/A _4592_/B vssd1 vssd1 vccd1 vccd1 _6393_/D sky130_fd_sc_hd__nor2_1
X_3543_ _3544_/A _3544_/B vssd1 vssd1 vccd1 vccd1 _3545_/B sky130_fd_sc_hd__nand2_1
X_3474_ _3474_/A vssd1 vssd1 vccd1 vccd1 _6315_/D sky130_fd_sc_hd__clkbuf_1
X_6262_ _6808_/Q _6247_/X _6261_/Y _6255_/X vssd1 vssd1 vccd1 vccd1 _6808_/D sky130_fd_sc_hd__o211a_1
XFILLER_103_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5213_ _5213_/A vssd1 vssd1 vccd1 vccd1 _6586_/D sky130_fd_sc_hd__clkbuf_1
X_6193_ _6787_/Q _5342_/X _6192_/X _6190_/X vssd1 vssd1 vccd1 vccd1 _6787_/D sky130_fd_sc_hd__o211a_1
X_5144_ _6692_/Q _6724_/Q _6756_/Q _6788_/Q _5126_/X _5138_/X vssd1 vssd1 vccd1 vccd1
+ _5144_/X sky130_fd_sc_hd__mux4_2
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5075_ _5118_/B vssd1 vssd1 vccd1 vccd1 _5075_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4026_ _4026_/A _4026_/B _4026_/C vssd1 vssd1 vccd1 vccd1 _4026_/X sky130_fd_sc_hd__and3_1
XFILLER_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6822__82 vssd1 vssd1 vccd1 vccd1 _6822__82/HI _6931_/A sky130_fd_sc_hd__conb_1
X_5977_ _6478_/Q _6056_/B _6056_/C _5976_/X vssd1 vssd1 vccd1 vccd1 _5977_/X sky130_fd_sc_hd__a31o_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4928_ _4928_/A _4928_/B vssd1 vssd1 vccd1 vccd1 _4928_/X sky130_fd_sc_hd__and2_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _5273_/A vssd1 vssd1 vccd1 vccd1 _4959_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6529_ _6554_/CLK _6529_/D vssd1 vssd1 vccd1 vccd1 _6529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _3193_/A vssd1 vssd1 vccd1 vccd1 _3190_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _6723_/Q _5888_/X _5899_/X _5863_/X vssd1 vssd1 vccd1 vccd1 _6723_/D sky130_fd_sc_hd__o211a_1
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5831_ _5602_/X _5830_/X _5842_/S vssd1 vssd1 vccd1 vccd1 _5831_/X sky130_fd_sc_hd__mux2_1
X_5762_ _6280_/A _5734_/X _5735_/X _5761_/X _5743_/X vssd1 vssd1 vccd1 vccd1 _5762_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4713_ _4735_/A vssd1 vssd1 vccd1 vccd1 _4722_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5693_ _5524_/X _5692_/X _5721_/S vssd1 vssd1 vccd1 vccd1 _5693_/X sky130_fd_sc_hd__mux2_1
X_4644_ _4644_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _4644_/X sky130_fd_sc_hd__or2_1
X_4575_ _4622_/A _4512_/B _4547_/B _4623_/A vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__a22oi_1
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6314_ _6531_/CLK _6314_/D vssd1 vssd1 vccd1 vccd1 _6314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3526_ _3526_/A _3539_/B _3524_/X vssd1 vssd1 vccd1 vccd1 _3544_/A sky130_fd_sc_hd__or3b_1
X_6245_ _6227_/X _6243_/Y _6244_/X vssd1 vssd1 vccd1 vccd1 _6245_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3457_ _3457_/A vssd1 vssd1 vccd1 vccd1 _6307_/D sky130_fd_sc_hd__clkbuf_1
X_3388_ _6291_/Q _3390_/C _3398_/B vssd1 vssd1 vccd1 vccd1 _3388_/Y sky130_fd_sc_hd__o21ai_1
X_6176_ _6780_/Q _6169_/X _6175_/X _6165_/X vssd1 vssd1 vccd1 vccd1 _6780_/D sky130_fd_sc_hd__o211a_1
X_5127_ _6689_/Q _6721_/Q _6753_/Q _6785_/Q _5126_/X _4950_/A vssd1 vssd1 vccd1 vccd1
+ _5127_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5058_ _6678_/Q _6710_/Q _6742_/Q _6774_/Q _5049_/X _5029_/X vssd1 vssd1 vccd1 vccd1
+ _5059_/B sky130_fd_sc_hd__mux4_1
XFILLER_84_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4009_ _4009_/A _4009_/B _4009_/C vssd1 vssd1 vccd1 vccd1 _4019_/B sky130_fd_sc_hd__nand3_2
XFILLER_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_3 _5570_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _6379_/Q vssd1 vssd1 vccd1 vccd1 _4547_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3311_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3311_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4291_ _4296_/A _4449_/A _4300_/B _4296_/C vssd1 vssd1 vccd1 vccd1 _4304_/A sky130_fd_sc_hd__nand4_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6030_ _6746_/Q _5619_/X _6044_/S vssd1 vssd1 vccd1 vccd1 _6030_/X sky130_fd_sc_hd__mux2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3242_ _3243_/A vssd1 vssd1 vccd1 vccd1 _3242_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6932_ _6932_/A _3227_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5814_ _5570_/X _5813_/X _5814_/S vssd1 vssd1 vccd1 vccd1 _5814_/X sky130_fd_sc_hd__mux2_1
X_6794_ _6795_/CLK _6794_/D vssd1 vssd1 vccd1 vccd1 _6794_/Q sky130_fd_sc_hd__dfxtp_1
X_5745_ _6697_/Q _5718_/X _5744_/X _5739_/X vssd1 vssd1 vccd1 vccd1 _6697_/D sky130_fd_sc_hd__o211a_1
X_5676_ _5880_/A _5880_/B vssd1 vssd1 vccd1 vccd1 _6062_/C sky130_fd_sc_hd__and2b_1
XFILLER_30_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4627_ _4627_/A _4627_/B vssd1 vssd1 vccd1 vccd1 _4642_/B sky130_fd_sc_hd__xnor2_2
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4558_ _4518_/B _4541_/Y _4572_/A _4557_/X vssd1 vssd1 vccd1 vccd1 _4573_/B sky130_fd_sc_hd__o211a_2
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4489_ _4545_/D vssd1 vssd1 vccd1 vccd1 _4597_/B sky130_fd_sc_hd__clkbuf_2
X_3509_ _6649_/Q vssd1 vssd1 vccd1 vccd1 _3661_/A sky130_fd_sc_hd__clkbuf_2
X_6228_ _6249_/A vssd1 vssd1 vccd1 vccd1 _6243_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6159_ _6773_/Q _6156_/X _6158_/X _6152_/X vssd1 vssd1 vccd1 vccd1 _6773_/D sky130_fd_sc_hd__o211a_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6842__102 vssd1 vssd1 vccd1 vccd1 _6842__102/HI _6951_/A sky130_fd_sc_hd__conb_1
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _3860_/A _3860_/B vssd1 vssd1 vccd1 vccd1 _6348_/D sky130_fd_sc_hd__nor2_1
X_3791_ _3810_/A _3792_/B _3792_/C vssd1 vssd1 vccd1 vccd1 _3793_/A sky130_fd_sc_hd__a21oi_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5530_ _6673_/Q _5529_/X _5562_/S vssd1 vssd1 vccd1 vccd1 _5531_/B sky130_fd_sc_hd__mux2_1
X_5461_ _5474_/A _5461_/B vssd1 vssd1 vccd1 vccd1 _5462_/A sky130_fd_sc_hd__and2_1
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4412_ _4428_/B _4428_/C _4428_/A vssd1 vssd1 vccd1 vccd1 _4414_/B sky130_fd_sc_hd__a21oi_1
X_5392_ _6638_/Q _5396_/B vssd1 vssd1 vccd1 vccd1 _5393_/A sky130_fd_sc_hd__and2_1
X_4343_ _4418_/A _4343_/B vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__and2_1
XFILLER_113_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4274_ _4274_/A vssd1 vssd1 vccd1 vccd1 _6380_/D sky130_fd_sc_hd__clkbuf_1
X_3225_ input1/X vssd1 vssd1 vccd1 vccd1 _3250_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6013_ _6040_/A vssd1 vssd1 vccd1 vccd1 _6013_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6915_ _6915_/A _3206_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__ebufn_8
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6777_ _6532_/Q _6777_/D vssd1 vssd1 vccd1 vccd1 _6777_/Q sky130_fd_sc_hd__dfxtp_1
X_3989_ _3986_/X _5239_/B _3989_/C vssd1 vssd1 vccd1 vccd1 _3990_/A sky130_fd_sc_hd__and3b_1
X_5728_ _6694_/Q _5380_/X _5726_/X _5727_/X _5707_/X vssd1 vssd1 vccd1 vccd1 _6694_/D
+ sky130_fd_sc_hd__o221a_1
X_5659_ _6476_/Q vssd1 vssd1 vccd1 vccd1 _5659_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _4935_/X _4936_/X _6543_/Q vssd1 vssd1 vccd1 vccd1 _4962_/B sky130_fd_sc_hd__a21oi_1
X_6700_ _6799_/CLK _6700_/D vssd1 vssd1 vccd1 vccd1 _6700_/Q sky130_fd_sc_hd__dfxtp_1
X_4892_ _6513_/Q _4887_/X _4888_/X input40/X vssd1 vssd1 vccd1 vccd1 _6513_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3912_ _3909_/Y _3911_/X _3913_/A vssd1 vssd1 vccd1 vccd1 _3914_/B sky130_fd_sc_hd__a21bo_1
X_6631_ _6799_/CLK _6631_/D vssd1 vssd1 vccd1 vccd1 _6631_/Q sky130_fd_sc_hd__dfxtp_1
X_3843_ _3843_/A _3843_/B vssd1 vssd1 vccd1 vccd1 _3843_/Y sky130_fd_sc_hd__xnor2_1
Xrepeater70 _6795_/CLK vssd1 vssd1 vccd1 vccd1 _6763_/CLK sky130_fd_sc_hd__buf_12
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3774_ _3741_/A _3741_/C _3741_/B vssd1 vssd1 vccd1 vccd1 _3775_/C sky130_fd_sc_hd__a21boi_1
X_6562_ _6562_/CLK _6562_/D vssd1 vssd1 vccd1 vccd1 _6900_/A sky130_fd_sc_hd__dfxtp_1
X_5513_ _5971_/A _6629_/Q _5971_/B vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__or3b_4
X_6493_ _6795_/CLK _6493_/D vssd1 vssd1 vccd1 vccd1 _6493_/Q sky130_fd_sc_hd__dfxtp_2
X_5444_ _5444_/A vssd1 vssd1 vccd1 vccd1 _6655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5375_ _6634_/Q _5396_/B vssd1 vssd1 vccd1 vccd1 _5376_/A sky130_fd_sc_hd__and2_1
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4326_ _4326_/A vssd1 vssd1 vccd1 vccd1 _6385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4257_ _4257_/A _4257_/B vssd1 vssd1 vccd1 vccd1 _4258_/A sky130_fd_sc_hd__and2_1
XFILLER_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3208_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3208_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4188_ _4188_/A vssd1 vssd1 vccd1 vccd1 _4188_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3490_ _3490_/A vssd1 vssd1 vccd1 vccd1 _6322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5160_ _5160_/A _5160_/B _5160_/C vssd1 vssd1 vccd1 vccd1 _5161_/A sky130_fd_sc_hd__and3_1
XFILLER_68_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5091_ _6683_/Q _6715_/Q _6747_/Q _6779_/Q _5083_/X _5063_/X vssd1 vssd1 vccd1 vccd1
+ _5092_/B sky130_fd_sc_hd__mux4_1
X_4111_ _4109_/X _4220_/A _3781_/X vssd1 vssd1 vccd1 vccd1 _4111_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4042_ _4042_/A _4042_/B _4042_/C vssd1 vssd1 vccd1 vccd1 _4043_/C sky130_fd_sc_hd__nand3_1
XFILLER_110_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _6739_/Q _5984_/X _5992_/X _5959_/X vssd1 vssd1 vccd1 vccd1 _6739_/D sky130_fd_sc_hd__o211a_1
XFILLER_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4944_ _5118_/B vssd1 vssd1 vccd1 vccd1 _5041_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4875_ _6501_/Q _4870_/X _4873_/X input47/X vssd1 vssd1 vccd1 vccd1 _6501_/D sky130_fd_sc_hd__a22o_1
X_6614_ _6667_/CLK _6614_/D vssd1 vssd1 vccd1 vccd1 _6614_/Q sky130_fd_sc_hd__dfxtp_1
X_3826_ _3826_/A _3826_/B vssd1 vssd1 vccd1 vccd1 _3826_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6545_ _6546_/CLK _6545_/D vssd1 vssd1 vccd1 vccd1 _6545_/Q sky130_fd_sc_hd__dfxtp_1
X_3757_ _3757_/A vssd1 vssd1 vccd1 vccd1 _3810_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6476_ _6763_/CLK _6476_/D vssd1 vssd1 vccd1 vccd1 _6476_/Q sky130_fd_sc_hd__dfxtp_1
X_3688_ _3729_/A _3755_/D vssd1 vssd1 vccd1 vccd1 _3692_/A sky130_fd_sc_hd__nand2_1
X_5427_ _5427_/A vssd1 vssd1 vccd1 vccd1 _6650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5358_ _6628_/Q vssd1 vssd1 vccd1 vccd1 _5882_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4309_ _4479_/B _6666_/Q _4433_/C _4400_/D vssd1 vssd1 vccd1 vccd1 _4354_/C sky130_fd_sc_hd__and4_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5289_ _5289_/A vssd1 vssd1 vccd1 vccd1 _6608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4660_ _6338_/Q _4666_/B vssd1 vssd1 vccd1 vccd1 _4661_/A sky130_fd_sc_hd__and2_1
X_3611_ _3611_/A _3648_/A vssd1 vssd1 vccd1 vccd1 _3641_/C sky130_fd_sc_hd__nor2_1
X_6330_ _6554_/CLK _6330_/D vssd1 vssd1 vccd1 vccd1 _6330_/Q sky130_fd_sc_hd__dfxtp_1
X_4591_ _4591_/A _4615_/D vssd1 vssd1 vccd1 vccd1 _4592_/B sky130_fd_sc_hd__xor2_1
X_3542_ _3565_/A _3542_/B vssd1 vssd1 vccd1 vccd1 _3544_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3473_ _6315_/Q _6519_/Q _3473_/S vssd1 vssd1 vccd1 vccd1 _3474_/A sky130_fd_sc_hd__mux2_1
X_6261_ _6248_/X _6260_/Y _6244_/X vssd1 vssd1 vccd1 vccd1 _6261_/Y sky130_fd_sc_hd__o21ai_1
X_5212_ _5243_/A _5212_/B _5212_/C vssd1 vssd1 vccd1 vccd1 _5213_/A sky130_fd_sc_hd__and3_1
XFILLER_88_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6192_ _6240_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _6192_/X sky130_fd_sc_hd__or2_1
X_5143_ _6913_/A _5149_/B vssd1 vssd1 vccd1 vccd1 _5147_/B sky130_fd_sc_hd__or2_1
XFILLER_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5074_ _6901_/A _5041_/X _5073_/X _5068_/X vssd1 vssd1 vccd1 vccd1 _6563_/D sky130_fd_sc_hd__o211a_1
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4025_ _3985_/A _3985_/B _4024_/Y vssd1 vssd1 vccd1 vccd1 _4026_/C sky130_fd_sc_hd__a21o_1
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5976_ _6003_/A vssd1 vssd1 vccd1 vccd1 _5976_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4927_ _4927_/A vssd1 vssd1 vccd1 vccd1 _6530_/D sky130_fd_sc_hd__clkbuf_1
X_4858_ _5284_/A vssd1 vssd1 vccd1 vccd1 _5273_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3809_ _3809_/A _3809_/B vssd1 vssd1 vccd1 vccd1 _3811_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4789_ _6412_/Q _4789_/B vssd1 vssd1 vccd1 vccd1 _4790_/A sky130_fd_sc_hd__and2_1
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6528_ _6528_/CLK _6528_/D vssd1 vssd1 vccd1 vccd1 _6528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6459_ _6789_/CLK _6459_/D vssd1 vssd1 vccd1 vccd1 _6459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5830_ _6712_/Q _5603_/X _5841_/S vssd1 vssd1 vccd1 vccd1 _5830_/X sky130_fd_sc_hd__mux2_1
X_5761_ _5651_/X _5760_/X _5771_/S vssd1 vssd1 vccd1 vccd1 _5761_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4712_ _4712_/A vssd1 vssd1 vccd1 vccd1 _6425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5692_ _6689_/Q _5529_/X _5764_/S vssd1 vssd1 vccd1 vccd1 _5692_/X sky130_fd_sc_hd__mux2_1
X_4643_ _4642_/A _4642_/B _4642_/C vssd1 vssd1 vccd1 vccd1 _4644_/B sky130_fd_sc_hd__a21oi_1
X_4574_ _4574_/A _4597_/B vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__nand2_1
X_6313_ _6528_/CLK _6313_/D vssd1 vssd1 vccd1 vccd1 _6313_/Q sky130_fd_sc_hd__dfxtp_1
X_3525_ _3522_/Y _3524_/X _3526_/A vssd1 vssd1 vccd1 vccd1 _3527_/B sky130_fd_sc_hd__a21bo_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _6264_/A vssd1 vssd1 vccd1 vccd1 _6244_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3456_ _6307_/Q _6511_/Q _3462_/S vssd1 vssd1 vccd1 vccd1 _3457_/A sky130_fd_sc_hd__mux2_1
X_3387_ _3392_/C vssd1 vssd1 vccd1 vccd1 _3398_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6175_ _6277_/A _6180_/B vssd1 vssd1 vccd1 vccd1 _6175_/X sky130_fd_sc_hd__or2_1
XFILLER_84_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5126_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5057_ _6898_/A _5041_/X _5056_/X _5034_/X vssd1 vssd1 vccd1 vccd1 _6560_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4008_ _4036_/A _4057_/B _4036_/C vssd1 vssd1 vccd1 vccd1 _4009_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5959_ _5999_/A vssd1 vssd1 vccd1 vccd1 _5959_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _3331_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3310_ _3310_/A vssd1 vssd1 vccd1 vccd1 _3310_/Y sky130_fd_sc_hd__inv_2
X_4290_ _4499_/A _4300_/B _4296_/C _4283_/A vssd1 vssd1 vccd1 vccd1 _4292_/B sky130_fd_sc_hd__a22o_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3243_/A vssd1 vssd1 vccd1 vccd1 _3241_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6931_ _6931_/A _3224_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5813_ _6709_/Q _5572_/X _5813_/S vssd1 vssd1 vccd1 vccd1 _5813_/X sky130_fd_sc_hd__mux2_1
X_6793_ _6795_/CLK _6793_/D vssd1 vssd1 vccd1 vccd1 _6793_/Q sky130_fd_sc_hd__dfxtp_1
X_5744_ _6263_/A _5734_/X _5735_/X _5742_/X _5743_/X vssd1 vssd1 vccd1 vccd1 _5744_/X
+ sky130_fd_sc_hd__a221o_1
X_5675_ _6478_/Q vssd1 vssd1 vccd1 vccd1 _6229_/A sky130_fd_sc_hd__buf_4
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4626_ _4626_/A _4626_/B vssd1 vssd1 vccd1 vccd1 _4627_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4557_ _4557_/A _4557_/B _4557_/C vssd1 vssd1 vccd1 vccd1 _4557_/X sky130_fd_sc_hd__or3_2
XFILLER_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4488_ _4442_/B _4487_/Y _4296_/A _4545_/D vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__o211a_1
X_3508_ _5162_/A vssd1 vssd1 vccd1 vccd1 _3899_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3439_ _3808_/C vssd1 vssd1 vccd1 vccd1 _5214_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6227_ _6248_/A vssd1 vssd1 vccd1 vccd1 _6227_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6158_ _6250_/A _6167_/B vssd1 vssd1 vccd1 vccd1 _6158_/X sky130_fd_sc_hd__or2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _6814_/Q _5109_/B vssd1 vssd1 vccd1 vccd1 _5109_/X sky130_fd_sc_hd__or2_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6756_/Q _6080_/X _6088_/X _6076_/X vssd1 vssd1 vccd1 vccd1 _6090_/B sky130_fd_sc_hd__a22o_1
XFILLER_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6881__141 vssd1 vssd1 vccd1 vccd1 _6881__141/HI _6990_/A sky130_fd_sc_hd__conb_1
XFILLER_76_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ _3790_/A _3813_/A vssd1 vssd1 vccd1 vccd1 _3792_/C sky130_fd_sc_hd__nor2_1
XFILLER_32_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5460_ _6308_/Q _4177_/A _5466_/S vssd1 vssd1 vccd1 vccd1 _5461_/B sky130_fd_sc_hd__mux2_1
X_4411_ _4427_/A _4411_/B vssd1 vssd1 vccd1 vccd1 _4428_/A sky130_fd_sc_hd__xnor2_1
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5391_ _5879_/A _5391_/B vssd1 vssd1 vccd1 vccd1 _6637_/D sky130_fd_sc_hd__nor2_1
X_4342_ _4342_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4343_/B sky130_fd_sc_hd__or2_1
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4273_ _4273_/A _4655_/B vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__and2_1
XFILLER_113_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6012_ _6743_/Q _5593_/X _6017_/S vssd1 vssd1 vccd1 vccd1 _6012_/X sky130_fd_sc_hd__mux2_1
X_3224_ _3224_/A vssd1 vssd1 vccd1 vccd1 _3224_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

