magic
tech sky130B
magscale 1 2
timestamp 1661702288
<< obsli1 >>
rect 1104 2159 68816 237745
<< obsm1 >>
rect 14 1912 69630 237776
<< metal2 >>
rect 1278 239200 1390 240000
rect 3854 239200 3966 240000
rect 6430 239200 6542 240000
rect 9006 239200 9118 240000
rect 12226 239200 12338 240000
rect 14802 239200 14914 240000
rect 17378 239200 17490 240000
rect 19954 239200 20066 240000
rect 22530 239200 22642 240000
rect 25750 239200 25862 240000
rect 28326 239200 28438 240000
rect 30902 239200 31014 240000
rect 33478 239200 33590 240000
rect 36054 239200 36166 240000
rect 38630 239200 38742 240000
rect 41850 239200 41962 240000
rect 44426 239200 44538 240000
rect 47002 239200 47114 240000
rect 49578 239200 49690 240000
rect 52154 239200 52266 240000
rect 55374 239200 55486 240000
rect 57950 239200 58062 240000
rect 60526 239200 60638 240000
rect 63102 239200 63214 240000
rect 65678 239200 65790 240000
rect 68254 239200 68366 240000
rect -10 0 102 800
rect 2566 0 2678 800
rect 5142 0 5254 800
rect 7718 0 7830 800
rect 10294 0 10406 800
rect 12870 0 12982 800
rect 16090 0 16202 800
rect 18666 0 18778 800
rect 21242 0 21354 800
rect 23818 0 23930 800
rect 26394 0 26506 800
rect 28970 0 29082 800
rect 32190 0 32302 800
rect 34766 0 34878 800
rect 37342 0 37454 800
rect 39918 0 40030 800
rect 42494 0 42606 800
rect 45714 0 45826 800
rect 48290 0 48402 800
rect 50866 0 50978 800
rect 53442 0 53554 800
rect 56018 0 56130 800
rect 58594 0 58706 800
rect 61814 0 61926 800
rect 64390 0 64502 800
rect 66966 0 67078 800
rect 69542 0 69654 800
<< obsm2 >>
rect 20 239144 1222 239442
rect 1446 239144 3798 239442
rect 4022 239144 6374 239442
rect 6598 239144 8950 239442
rect 9174 239144 12170 239442
rect 12394 239144 14746 239442
rect 14970 239144 17322 239442
rect 17546 239144 19898 239442
rect 20122 239144 22474 239442
rect 22698 239144 25694 239442
rect 25918 239144 28270 239442
rect 28494 239144 30846 239442
rect 31070 239144 33422 239442
rect 33646 239144 35998 239442
rect 36222 239144 38574 239442
rect 38798 239144 41794 239442
rect 42018 239144 44370 239442
rect 44594 239144 46946 239442
rect 47170 239144 49522 239442
rect 49746 239144 52098 239442
rect 52322 239144 55318 239442
rect 55542 239144 57894 239442
rect 58118 239144 60470 239442
rect 60694 239144 63046 239442
rect 63270 239144 65622 239442
rect 65846 239144 68198 239442
rect 68422 239144 69624 239442
rect 20 856 69624 239144
rect 158 734 2510 856
rect 2734 734 5086 856
rect 5310 734 7662 856
rect 7886 734 10238 856
rect 10462 734 12814 856
rect 13038 734 16034 856
rect 16258 734 18610 856
rect 18834 734 21186 856
rect 21410 734 23762 856
rect 23986 734 26338 856
rect 26562 734 28914 856
rect 29138 734 32134 856
rect 32358 734 34710 856
rect 34934 734 37286 856
rect 37510 734 39862 856
rect 40086 734 42438 856
rect 42662 734 45658 856
rect 45882 734 48234 856
rect 48458 734 50810 856
rect 51034 734 53386 856
rect 53610 734 55962 856
rect 56186 734 58538 856
rect 58762 734 61758 856
rect 61982 734 64334 856
rect 64558 734 66910 856
rect 67134 734 69486 856
<< metal3 >>
rect 0 238628 800 238868
rect 69200 237948 70000 238188
rect 0 235908 800 236148
rect 69200 235228 70000 235468
rect 0 232508 800 232748
rect 69200 232508 70000 232748
rect 0 229788 800 230028
rect 69200 229788 70000 230028
rect 0 227068 800 227308
rect 69200 227068 70000 227308
rect 0 224348 800 224588
rect 69200 224348 70000 224588
rect 0 221628 800 221868
rect 69200 220948 70000 221188
rect 0 218228 800 218468
rect 69200 218228 70000 218468
rect 0 215508 800 215748
rect 69200 215508 70000 215748
rect 0 212788 800 213028
rect 69200 212788 70000 213028
rect 0 210068 800 210308
rect 69200 210068 70000 210308
rect 0 207348 800 207588
rect 69200 206668 70000 206908
rect 0 204628 800 204868
rect 69200 203948 70000 204188
rect 0 201228 800 201468
rect 69200 201228 70000 201468
rect 0 198508 800 198748
rect 69200 198508 70000 198748
rect 0 195788 800 196028
rect 69200 195788 70000 196028
rect 0 193068 800 193308
rect 69200 193068 70000 193308
rect 0 190348 800 190588
rect 69200 189668 70000 189908
rect 0 186948 800 187188
rect 69200 186948 70000 187188
rect 0 184228 800 184468
rect 69200 184228 70000 184468
rect 0 181508 800 181748
rect 69200 181508 70000 181748
rect 0 178788 800 179028
rect 69200 178788 70000 179028
rect 0 176068 800 176308
rect 69200 175388 70000 175628
rect 0 173348 800 173588
rect 69200 172668 70000 172908
rect 0 169948 800 170188
rect 69200 169948 70000 170188
rect 0 167228 800 167468
rect 69200 167228 70000 167468
rect 0 164508 800 164748
rect 69200 164508 70000 164748
rect 0 161788 800 162028
rect 69200 161788 70000 162028
rect 0 159068 800 159308
rect 69200 158388 70000 158628
rect 0 155668 800 155908
rect 69200 155668 70000 155908
rect 0 152948 800 153188
rect 69200 152948 70000 153188
rect 0 150228 800 150468
rect 69200 150228 70000 150468
rect 0 147508 800 147748
rect 69200 147508 70000 147748
rect 0 144788 800 145028
rect 69200 144108 70000 144348
rect 0 142068 800 142308
rect 69200 141388 70000 141628
rect 0 138668 800 138908
rect 69200 138668 70000 138908
rect 0 135948 800 136188
rect 69200 135948 70000 136188
rect 0 133228 800 133468
rect 69200 133228 70000 133468
rect 0 130508 800 130748
rect 69200 130508 70000 130748
rect 0 127788 800 128028
rect 69200 127108 70000 127348
rect 0 124388 800 124628
rect 69200 124388 70000 124628
rect 0 121668 800 121908
rect 69200 121668 70000 121908
rect 0 118948 800 119188
rect 69200 118948 70000 119188
rect 0 116228 800 116468
rect 69200 116228 70000 116468
rect 0 113508 800 113748
rect 69200 112828 70000 113068
rect 0 110788 800 111028
rect 69200 110108 70000 110348
rect 0 107388 800 107628
rect 69200 107388 70000 107628
rect 0 104668 800 104908
rect 69200 104668 70000 104908
rect 0 101948 800 102188
rect 69200 101948 70000 102188
rect 0 99228 800 99468
rect 69200 99228 70000 99468
rect 0 96508 800 96748
rect 69200 95828 70000 96068
rect 0 93108 800 93348
rect 69200 93108 70000 93348
rect 0 90388 800 90628
rect 69200 90388 70000 90628
rect 0 87668 800 87908
rect 69200 87668 70000 87908
rect 0 84948 800 85188
rect 69200 84948 70000 85188
rect 0 82228 800 82468
rect 69200 81548 70000 81788
rect 0 79508 800 79748
rect 69200 78828 70000 79068
rect 0 76108 800 76348
rect 69200 76108 70000 76348
rect 0 73388 800 73628
rect 69200 73388 70000 73628
rect 0 70668 800 70908
rect 69200 70668 70000 70908
rect 0 67948 800 68188
rect 69200 67948 70000 68188
rect 0 65228 800 65468
rect 69200 64548 70000 64788
rect 0 61828 800 62068
rect 69200 61828 70000 62068
rect 0 59108 800 59348
rect 69200 59108 70000 59348
rect 0 56388 800 56628
rect 69200 56388 70000 56628
rect 0 53668 800 53908
rect 69200 53668 70000 53908
rect 0 50948 800 51188
rect 69200 50268 70000 50508
rect 0 48228 800 48468
rect 69200 47548 70000 47788
rect 0 44828 800 45068
rect 69200 44828 70000 45068
rect 0 42108 800 42348
rect 69200 42108 70000 42348
rect 0 39388 800 39628
rect 69200 39388 70000 39628
rect 0 36668 800 36908
rect 69200 36668 70000 36908
rect 0 33948 800 34188
rect 69200 33268 70000 33508
rect 0 30548 800 30788
rect 69200 30548 70000 30788
rect 0 27828 800 28068
rect 69200 27828 70000 28068
rect 0 25108 800 25348
rect 69200 25108 70000 25348
rect 0 22388 800 22628
rect 69200 22388 70000 22628
rect 0 19668 800 19908
rect 69200 18988 70000 19228
rect 0 16948 800 17188
rect 69200 16268 70000 16508
rect 0 13548 800 13788
rect 69200 13548 70000 13788
rect 0 10828 800 11068
rect 69200 10828 70000 11068
rect 0 8108 800 8348
rect 69200 8108 70000 8348
rect 0 5388 800 5628
rect 69200 5388 70000 5628
rect 0 2668 800 2908
rect 69200 1988 70000 2228
<< obsm3 >>
rect 880 238548 69306 238781
rect 800 238268 69306 238548
rect 800 237868 69120 238268
rect 800 236228 69306 237868
rect 880 235828 69306 236228
rect 800 235548 69306 235828
rect 800 235148 69120 235548
rect 800 232828 69306 235148
rect 880 232428 69120 232828
rect 800 230108 69306 232428
rect 880 229708 69120 230108
rect 800 227388 69306 229708
rect 880 226988 69120 227388
rect 800 224668 69306 226988
rect 880 224268 69120 224668
rect 800 221948 69306 224268
rect 880 221548 69306 221948
rect 800 221268 69306 221548
rect 800 220868 69120 221268
rect 800 218548 69306 220868
rect 880 218148 69120 218548
rect 800 215828 69306 218148
rect 880 215428 69120 215828
rect 800 213108 69306 215428
rect 880 212708 69120 213108
rect 800 210388 69306 212708
rect 880 209988 69120 210388
rect 800 207668 69306 209988
rect 880 207268 69306 207668
rect 800 206988 69306 207268
rect 800 206588 69120 206988
rect 800 204948 69306 206588
rect 880 204548 69306 204948
rect 800 204268 69306 204548
rect 800 203868 69120 204268
rect 800 201548 69306 203868
rect 880 201148 69120 201548
rect 800 198828 69306 201148
rect 880 198428 69120 198828
rect 800 196108 69306 198428
rect 880 195708 69120 196108
rect 800 193388 69306 195708
rect 880 192988 69120 193388
rect 800 190668 69306 192988
rect 880 190268 69306 190668
rect 800 189988 69306 190268
rect 800 189588 69120 189988
rect 800 187268 69306 189588
rect 880 186868 69120 187268
rect 800 184548 69306 186868
rect 880 184148 69120 184548
rect 800 181828 69306 184148
rect 880 181428 69120 181828
rect 800 179108 69306 181428
rect 880 178708 69120 179108
rect 800 176388 69306 178708
rect 880 175988 69306 176388
rect 800 175708 69306 175988
rect 800 175308 69120 175708
rect 800 173668 69306 175308
rect 880 173268 69306 173668
rect 800 172988 69306 173268
rect 800 172588 69120 172988
rect 800 170268 69306 172588
rect 880 169868 69120 170268
rect 800 167548 69306 169868
rect 880 167148 69120 167548
rect 800 164828 69306 167148
rect 880 164428 69120 164828
rect 800 162108 69306 164428
rect 880 161708 69120 162108
rect 800 159388 69306 161708
rect 880 158988 69306 159388
rect 800 158708 69306 158988
rect 800 158308 69120 158708
rect 800 155988 69306 158308
rect 880 155588 69120 155988
rect 800 153268 69306 155588
rect 880 152868 69120 153268
rect 800 150548 69306 152868
rect 880 150148 69120 150548
rect 800 147828 69306 150148
rect 880 147428 69120 147828
rect 800 145108 69306 147428
rect 880 144708 69306 145108
rect 800 144428 69306 144708
rect 800 144028 69120 144428
rect 800 142388 69306 144028
rect 880 141988 69306 142388
rect 800 141708 69306 141988
rect 800 141308 69120 141708
rect 800 138988 69306 141308
rect 880 138588 69120 138988
rect 800 136268 69306 138588
rect 880 135868 69120 136268
rect 800 133548 69306 135868
rect 880 133148 69120 133548
rect 800 130828 69306 133148
rect 880 130428 69120 130828
rect 800 128108 69306 130428
rect 880 127708 69306 128108
rect 800 127428 69306 127708
rect 800 127028 69120 127428
rect 800 124708 69306 127028
rect 880 124308 69120 124708
rect 800 121988 69306 124308
rect 880 121588 69120 121988
rect 800 119268 69306 121588
rect 880 118868 69120 119268
rect 800 116548 69306 118868
rect 880 116148 69120 116548
rect 800 113828 69306 116148
rect 880 113428 69306 113828
rect 800 113148 69306 113428
rect 800 112748 69120 113148
rect 800 111108 69306 112748
rect 880 110708 69306 111108
rect 800 110428 69306 110708
rect 800 110028 69120 110428
rect 800 107708 69306 110028
rect 880 107308 69120 107708
rect 800 104988 69306 107308
rect 880 104588 69120 104988
rect 800 102268 69306 104588
rect 880 101868 69120 102268
rect 800 99548 69306 101868
rect 880 99148 69120 99548
rect 800 96828 69306 99148
rect 880 96428 69306 96828
rect 800 96148 69306 96428
rect 800 95748 69120 96148
rect 800 93428 69306 95748
rect 880 93028 69120 93428
rect 800 90708 69306 93028
rect 880 90308 69120 90708
rect 800 87988 69306 90308
rect 880 87588 69120 87988
rect 800 85268 69306 87588
rect 880 84868 69120 85268
rect 800 82548 69306 84868
rect 880 82148 69306 82548
rect 800 81868 69306 82148
rect 800 81468 69120 81868
rect 800 79828 69306 81468
rect 880 79428 69306 79828
rect 800 79148 69306 79428
rect 800 78748 69120 79148
rect 800 76428 69306 78748
rect 880 76028 69120 76428
rect 800 73708 69306 76028
rect 880 73308 69120 73708
rect 800 70988 69306 73308
rect 880 70588 69120 70988
rect 800 68268 69306 70588
rect 880 67868 69120 68268
rect 800 65548 69306 67868
rect 880 65148 69306 65548
rect 800 64868 69306 65148
rect 800 64468 69120 64868
rect 800 62148 69306 64468
rect 880 61748 69120 62148
rect 800 59428 69306 61748
rect 880 59028 69120 59428
rect 800 56708 69306 59028
rect 880 56308 69120 56708
rect 800 53988 69306 56308
rect 880 53588 69120 53988
rect 800 51268 69306 53588
rect 880 50868 69306 51268
rect 800 50588 69306 50868
rect 800 50188 69120 50588
rect 800 48548 69306 50188
rect 880 48148 69306 48548
rect 800 47868 69306 48148
rect 800 47468 69120 47868
rect 800 45148 69306 47468
rect 880 44748 69120 45148
rect 800 42428 69306 44748
rect 880 42028 69120 42428
rect 800 39708 69306 42028
rect 880 39308 69120 39708
rect 800 36988 69306 39308
rect 880 36588 69120 36988
rect 800 34268 69306 36588
rect 880 33868 69306 34268
rect 800 33588 69306 33868
rect 800 33188 69120 33588
rect 800 30868 69306 33188
rect 880 30468 69120 30868
rect 800 28148 69306 30468
rect 880 27748 69120 28148
rect 800 25428 69306 27748
rect 880 25028 69120 25428
rect 800 22708 69306 25028
rect 880 22308 69120 22708
rect 800 19988 69306 22308
rect 880 19588 69306 19988
rect 800 19308 69306 19588
rect 800 18908 69120 19308
rect 800 17268 69306 18908
rect 880 16868 69306 17268
rect 800 16588 69306 16868
rect 800 16188 69120 16588
rect 800 13868 69306 16188
rect 880 13468 69120 13868
rect 800 11148 69306 13468
rect 880 10748 69120 11148
rect 800 8428 69306 10748
rect 880 8028 69120 8428
rect 800 5708 69306 8028
rect 880 5308 69120 5708
rect 800 2988 69306 5308
rect 880 2588 69306 2988
rect 800 2308 69306 2588
rect 800 2075 69120 2308
<< metal4 >>
rect 4208 2128 4528 237776
rect 19568 2128 19888 237776
rect 34928 2128 35248 237776
rect 50288 2128 50608 237776
rect 65648 2128 65968 237776
<< obsm4 >>
rect 19379 3435 19488 228037
rect 19968 3435 34848 228037
rect 35328 3435 50208 228037
rect 50688 3435 55877 228037
<< labels >>
rlabel metal3 s 0 152948 800 153188 6 active
port 1 nsew signal input
rlabel metal3 s 69200 133228 70000 133468 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 69200 44828 70000 45068 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 69200 50268 70000 50508 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 io_in[12]
port 5 nsew signal input
rlabel metal3 s 69200 110108 70000 110348 6 io_in[13]
port 6 nsew signal input
rlabel metal3 s 69200 104668 70000 104908 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 56018 0 56130 800 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 69200 164508 70000 164748 6 io_in[17]
port 10 nsew signal input
rlabel metal3 s 69200 144108 70000 144348 6 io_in[18]
port 11 nsew signal input
rlabel metal3 s 69200 56388 70000 56628 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 204628 800 204868 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 69200 90388 70000 90628 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 69200 198508 70000 198748 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 0 176068 800 176308 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 47002 239200 47114 240000 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 0 104668 800 104908 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 57950 239200 58062 240000 6 io_in[25]
port 19 nsew signal input
rlabel metal3 s 0 229788 800 230028 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 69200 47548 70000 47788 6 io_in[27]
port 21 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 io_in[28]
port 22 nsew signal input
rlabel metal3 s 69200 30548 70000 30788 6 io_in[29]
port 23 nsew signal input
rlabel metal3 s 0 184228 800 184468 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 0 159068 800 159308 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 195788 800 196028 6 io_in[31]
port 26 nsew signal input
rlabel metal3 s 0 61828 800 62068 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 69200 93108 70000 93348 6 io_in[33]
port 28 nsew signal input
rlabel metal3 s 69200 10828 70000 11068 6 io_in[34]
port 29 nsew signal input
rlabel metal3 s 69200 138668 70000 138908 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 0 138668 800 138908 6 io_in[36]
port 31 nsew signal input
rlabel metal3 s 69200 189668 70000 189908 6 io_in[37]
port 32 nsew signal input
rlabel metal3 s 69200 61828 70000 62068 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 0 124388 800 124628 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 50866 0 50978 800 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 66966 0 67078 800 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 69200 59108 70000 59348 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 0 13548 800 13788 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 69200 33268 70000 33508 6 io_oeb[0]
port 40 nsew signal bidirectional
rlabel metal2 s 28326 239200 28438 240000 6 io_oeb[10]
port 41 nsew signal bidirectional
rlabel metal3 s 69200 67948 70000 68188 6 io_oeb[11]
port 42 nsew signal bidirectional
rlabel metal2 s 33478 239200 33590 240000 6 io_oeb[12]
port 43 nsew signal bidirectional
rlabel metal3 s 69200 178788 70000 179028 6 io_oeb[13]
port 44 nsew signal bidirectional
rlabel metal3 s 69200 210068 70000 210308 6 io_oeb[14]
port 45 nsew signal bidirectional
rlabel metal3 s 69200 175388 70000 175628 6 io_oeb[15]
port 46 nsew signal bidirectional
rlabel metal3 s 0 50948 800 51188 6 io_oeb[16]
port 47 nsew signal bidirectional
rlabel metal3 s 69200 5388 70000 5628 6 io_oeb[17]
port 48 nsew signal bidirectional
rlabel metal2 s 55374 239200 55486 240000 6 io_oeb[18]
port 49 nsew signal bidirectional
rlabel metal3 s 0 27828 800 28068 6 io_oeb[19]
port 50 nsew signal bidirectional
rlabel metal3 s 69200 95828 70000 96068 6 io_oeb[1]
port 51 nsew signal bidirectional
rlabel metal3 s 0 2668 800 2908 6 io_oeb[20]
port 52 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 io_oeb[21]
port 53 nsew signal bidirectional
rlabel metal3 s 69200 227068 70000 227308 6 io_oeb[22]
port 54 nsew signal bidirectional
rlabel metal2 s 41850 239200 41962 240000 6 io_oeb[23]
port 55 nsew signal bidirectional
rlabel metal2 s 12870 0 12982 800 6 io_oeb[24]
port 56 nsew signal bidirectional
rlabel metal2 s 48290 0 48402 800 6 io_oeb[25]
port 57 nsew signal bidirectional
rlabel metal3 s 69200 172668 70000 172908 6 io_oeb[26]
port 58 nsew signal bidirectional
rlabel metal3 s 69200 27828 70000 28068 6 io_oeb[27]
port 59 nsew signal bidirectional
rlabel metal3 s 0 48228 800 48468 6 io_oeb[28]
port 60 nsew signal bidirectional
rlabel metal3 s 0 227068 800 227308 6 io_oeb[29]
port 61 nsew signal bidirectional
rlabel metal3 s 0 113508 800 113748 6 io_oeb[2]
port 62 nsew signal bidirectional
rlabel metal3 s 0 167228 800 167468 6 io_oeb[30]
port 63 nsew signal bidirectional
rlabel metal2 s 65678 239200 65790 240000 6 io_oeb[31]
port 64 nsew signal bidirectional
rlabel metal2 s 3854 239200 3966 240000 6 io_oeb[32]
port 65 nsew signal bidirectional
rlabel metal3 s 69200 218228 70000 218468 6 io_oeb[33]
port 66 nsew signal bidirectional
rlabel metal3 s 69200 220948 70000 221188 6 io_oeb[34]
port 67 nsew signal bidirectional
rlabel metal3 s 0 76108 800 76348 6 io_oeb[35]
port 68 nsew signal bidirectional
rlabel metal2 s 44426 239200 44538 240000 6 io_oeb[36]
port 69 nsew signal bidirectional
rlabel metal3 s 69200 184228 70000 184468 6 io_oeb[37]
port 70 nsew signal bidirectional
rlabel metal3 s 0 181508 800 181748 6 io_oeb[3]
port 71 nsew signal bidirectional
rlabel metal3 s 69200 130508 70000 130748 6 io_oeb[4]
port 72 nsew signal bidirectional
rlabel metal3 s 0 127788 800 128028 6 io_oeb[5]
port 73 nsew signal bidirectional
rlabel metal3 s 0 169948 800 170188 6 io_oeb[6]
port 74 nsew signal bidirectional
rlabel metal3 s 69200 229788 70000 230028 6 io_oeb[7]
port 75 nsew signal bidirectional
rlabel metal3 s 69200 161788 70000 162028 6 io_oeb[8]
port 76 nsew signal bidirectional
rlabel metal3 s 0 65228 800 65468 6 io_oeb[9]
port 77 nsew signal bidirectional
rlabel metal3 s 0 144788 800 145028 6 io_out[0]
port 78 nsew signal bidirectional
rlabel metal3 s 0 5388 800 5628 6 io_out[10]
port 79 nsew signal bidirectional
rlabel metal3 s 69200 13548 70000 13788 6 io_out[11]
port 80 nsew signal bidirectional
rlabel metal3 s 0 67948 800 68188 6 io_out[12]
port 81 nsew signal bidirectional
rlabel metal2 s 12226 239200 12338 240000 6 io_out[13]
port 82 nsew signal bidirectional
rlabel metal2 s 68254 239200 68366 240000 6 io_out[14]
port 83 nsew signal bidirectional
rlabel metal3 s 0 101948 800 102188 6 io_out[15]
port 84 nsew signal bidirectional
rlabel metal2 s 16090 0 16202 800 6 io_out[16]
port 85 nsew signal bidirectional
rlabel metal3 s 0 212788 800 213028 6 io_out[17]
port 86 nsew signal bidirectional
rlabel metal3 s 69200 121668 70000 121908 6 io_out[18]
port 87 nsew signal bidirectional
rlabel metal2 s 49578 239200 49690 240000 6 io_out[19]
port 88 nsew signal bidirectional
rlabel metal3 s 0 8108 800 8348 6 io_out[1]
port 89 nsew signal bidirectional
rlabel metal3 s 0 56388 800 56628 6 io_out[20]
port 90 nsew signal bidirectional
rlabel metal3 s 69200 64548 70000 64788 6 io_out[21]
port 91 nsew signal bidirectional
rlabel metal2 s 63102 239200 63214 240000 6 io_out[22]
port 92 nsew signal bidirectional
rlabel metal2 s 19954 239200 20066 240000 6 io_out[23]
port 93 nsew signal bidirectional
rlabel metal3 s 69200 181508 70000 181748 6 io_out[24]
port 94 nsew signal bidirectional
rlabel metal3 s 0 116228 800 116468 6 io_out[25]
port 95 nsew signal bidirectional
rlabel metal3 s 69200 84948 70000 85188 6 io_out[26]
port 96 nsew signal bidirectional
rlabel metal3 s 69200 152948 70000 153188 6 io_out[27]
port 97 nsew signal bidirectional
rlabel metal2 s 9006 239200 9118 240000 6 io_out[28]
port 98 nsew signal bidirectional
rlabel metal2 s 30902 239200 31014 240000 6 io_out[29]
port 99 nsew signal bidirectional
rlabel metal3 s 69200 135948 70000 136188 6 io_out[2]
port 100 nsew signal bidirectional
rlabel metal3 s 0 10828 800 11068 6 io_out[30]
port 101 nsew signal bidirectional
rlabel metal2 s 17378 239200 17490 240000 6 io_out[31]
port 102 nsew signal bidirectional
rlabel metal3 s 0 193068 800 193308 6 io_out[32]
port 103 nsew signal bidirectional
rlabel metal3 s 0 218228 800 218468 6 io_out[33]
port 104 nsew signal bidirectional
rlabel metal2 s 1278 239200 1390 240000 6 io_out[34]
port 105 nsew signal bidirectional
rlabel metal3 s 69200 81548 70000 81788 6 io_out[35]
port 106 nsew signal bidirectional
rlabel metal3 s 0 33948 800 34188 6 io_out[36]
port 107 nsew signal bidirectional
rlabel metal3 s 69200 99228 70000 99468 6 io_out[37]
port 108 nsew signal bidirectional
rlabel metal2 s 23818 0 23930 800 6 io_out[3]
port 109 nsew signal bidirectional
rlabel metal3 s 0 84948 800 85188 6 io_out[4]
port 110 nsew signal bidirectional
rlabel metal3 s 0 238628 800 238868 6 io_out[5]
port 111 nsew signal bidirectional
rlabel metal3 s 69200 155668 70000 155908 6 io_out[6]
port 112 nsew signal bidirectional
rlabel metal3 s 69200 116228 70000 116468 6 io_out[7]
port 113 nsew signal bidirectional
rlabel metal3 s 0 147508 800 147748 6 io_out[8]
port 114 nsew signal bidirectional
rlabel metal3 s 69200 215508 70000 215748 6 io_out[9]
port 115 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 237776 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 237776 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 237776 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 237776 6 vssd1
port 117 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 237776 6 vssd1
port 117 nsew ground bidirectional
rlabel metal3 s 0 207348 800 207588 6 wb_clk_i
port 118 nsew signal input
rlabel metal3 s 69200 235228 70000 235468 6 wb_rst_i
port 119 nsew signal input
rlabel metal3 s 0 110788 800 111028 6 wbs_ack_o
port 120 nsew signal bidirectional
rlabel metal3 s 69200 186948 70000 187188 6 wbs_adr_i[0]
port 121 nsew signal input
rlabel metal3 s 69200 212788 70000 213028 6 wbs_adr_i[10]
port 122 nsew signal input
rlabel metal3 s 0 90388 800 90628 6 wbs_adr_i[11]
port 123 nsew signal input
rlabel metal2 s 7718 0 7830 800 6 wbs_adr_i[12]
port 124 nsew signal input
rlabel metal2 s 58594 0 58706 800 6 wbs_adr_i[13]
port 125 nsew signal input
rlabel metal3 s 69200 124388 70000 124628 6 wbs_adr_i[14]
port 126 nsew signal input
rlabel metal3 s 0 235908 800 236148 6 wbs_adr_i[15]
port 127 nsew signal input
rlabel metal2 s 69542 0 69654 800 6 wbs_adr_i[16]
port 128 nsew signal input
rlabel metal3 s 69200 112828 70000 113068 6 wbs_adr_i[17]
port 129 nsew signal input
rlabel metal3 s 69200 78828 70000 79068 6 wbs_adr_i[18]
port 130 nsew signal input
rlabel metal3 s 0 135948 800 136188 6 wbs_adr_i[19]
port 131 nsew signal input
rlabel metal3 s 0 99228 800 99468 6 wbs_adr_i[1]
port 132 nsew signal input
rlabel metal3 s 69200 169948 70000 170188 6 wbs_adr_i[20]
port 133 nsew signal input
rlabel metal3 s 0 121668 800 121908 6 wbs_adr_i[21]
port 134 nsew signal input
rlabel metal3 s 0 53668 800 53908 6 wbs_adr_i[22]
port 135 nsew signal input
rlabel metal3 s 69200 73388 70000 73628 6 wbs_adr_i[23]
port 136 nsew signal input
rlabel metal3 s 0 201228 800 201468 6 wbs_adr_i[24]
port 137 nsew signal input
rlabel metal2 s 61814 0 61926 800 6 wbs_adr_i[25]
port 138 nsew signal input
rlabel metal3 s 0 73388 800 73628 6 wbs_adr_i[26]
port 139 nsew signal input
rlabel metal3 s 0 96508 800 96748 6 wbs_adr_i[27]
port 140 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 wbs_adr_i[28]
port 141 nsew signal input
rlabel metal3 s 0 198508 800 198748 6 wbs_adr_i[29]
port 142 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 wbs_adr_i[2]
port 143 nsew signal input
rlabel metal3 s 0 173348 800 173588 6 wbs_adr_i[30]
port 144 nsew signal input
rlabel metal3 s 69200 101948 70000 102188 6 wbs_adr_i[31]
port 145 nsew signal input
rlabel metal3 s 69200 22388 70000 22628 6 wbs_adr_i[3]
port 146 nsew signal input
rlabel metal3 s 69200 206668 70000 206908 6 wbs_adr_i[4]
port 147 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 wbs_adr_i[5]
port 148 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 wbs_adr_i[6]
port 149 nsew signal input
rlabel metal3 s 0 186948 800 187188 6 wbs_adr_i[7]
port 150 nsew signal input
rlabel metal3 s 69200 53668 70000 53908 6 wbs_adr_i[8]
port 151 nsew signal input
rlabel metal3 s 0 93108 800 93348 6 wbs_adr_i[9]
port 152 nsew signal input
rlabel metal2 s 38630 239200 38742 240000 6 wbs_cyc_i
port 153 nsew signal input
rlabel metal3 s 0 155668 800 155908 6 wbs_dat_i[0]
port 154 nsew signal input
rlabel metal3 s 0 190348 800 190588 6 wbs_dat_i[10]
port 155 nsew signal input
rlabel metal3 s 0 215508 800 215748 6 wbs_dat_i[11]
port 156 nsew signal input
rlabel metal3 s 0 210068 800 210308 6 wbs_dat_i[12]
port 157 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 wbs_dat_i[13]
port 158 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 wbs_dat_i[14]
port 159 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 wbs_dat_i[15]
port 160 nsew signal input
rlabel metal3 s 69200 1988 70000 2228 6 wbs_dat_i[16]
port 161 nsew signal input
rlabel metal3 s 69200 232508 70000 232748 6 wbs_dat_i[17]
port 162 nsew signal input
rlabel metal3 s 0 161788 800 162028 6 wbs_dat_i[18]
port 163 nsew signal input
rlabel metal3 s 0 232508 800 232748 6 wbs_dat_i[19]
port 164 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 wbs_dat_i[1]
port 165 nsew signal input
rlabel metal3 s 69200 141388 70000 141628 6 wbs_dat_i[20]
port 166 nsew signal input
rlabel metal3 s 69200 201228 70000 201468 6 wbs_dat_i[21]
port 167 nsew signal input
rlabel metal3 s 0 70668 800 70908 6 wbs_dat_i[22]
port 168 nsew signal input
rlabel metal3 s 69200 167228 70000 167468 6 wbs_dat_i[23]
port 169 nsew signal input
rlabel metal3 s 0 133228 800 133468 6 wbs_dat_i[24]
port 170 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 wbs_dat_i[25]
port 171 nsew signal input
rlabel metal3 s 69200 224348 70000 224588 6 wbs_dat_i[26]
port 172 nsew signal input
rlabel metal2 s 6430 239200 6542 240000 6 wbs_dat_i[27]
port 173 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 wbs_dat_i[28]
port 174 nsew signal input
rlabel metal3 s 69200 147508 70000 147748 6 wbs_dat_i[29]
port 175 nsew signal input
rlabel metal3 s 69200 39388 70000 39628 6 wbs_dat_i[2]
port 176 nsew signal input
rlabel metal3 s 69200 107388 70000 107628 6 wbs_dat_i[30]
port 177 nsew signal input
rlabel metal3 s 0 142068 800 142308 6 wbs_dat_i[31]
port 178 nsew signal input
rlabel metal3 s 69200 70668 70000 70908 6 wbs_dat_i[3]
port 179 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 wbs_dat_i[4]
port 180 nsew signal input
rlabel metal2 s 64390 0 64502 800 6 wbs_dat_i[5]
port 181 nsew signal input
rlabel metal3 s 69200 127108 70000 127348 6 wbs_dat_i[6]
port 182 nsew signal input
rlabel metal3 s 69200 237948 70000 238188 6 wbs_dat_i[7]
port 183 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 wbs_dat_i[8]
port 184 nsew signal input
rlabel metal3 s 69200 76108 70000 76348 6 wbs_dat_i[9]
port 185 nsew signal input
rlabel metal3 s 0 59108 800 59348 6 wbs_dat_o[0]
port 186 nsew signal bidirectional
rlabel metal3 s 69200 150228 70000 150468 6 wbs_dat_o[10]
port 187 nsew signal bidirectional
rlabel metal2 s 2566 0 2678 800 6 wbs_dat_o[11]
port 188 nsew signal bidirectional
rlabel metal3 s 69200 203948 70000 204188 6 wbs_dat_o[12]
port 189 nsew signal bidirectional
rlabel metal2 s 60526 239200 60638 240000 6 wbs_dat_o[13]
port 190 nsew signal bidirectional
rlabel metal3 s 69200 87668 70000 87908 6 wbs_dat_o[14]
port 191 nsew signal bidirectional
rlabel metal2 s 52154 239200 52266 240000 6 wbs_dat_o[15]
port 192 nsew signal bidirectional
rlabel metal3 s 0 82228 800 82468 6 wbs_dat_o[16]
port 193 nsew signal bidirectional
rlabel metal3 s 0 87668 800 87908 6 wbs_dat_o[17]
port 194 nsew signal bidirectional
rlabel metal3 s 69200 25108 70000 25348 6 wbs_dat_o[18]
port 195 nsew signal bidirectional
rlabel metal2 s -10 0 102 800 6 wbs_dat_o[19]
port 196 nsew signal bidirectional
rlabel metal3 s 69200 42108 70000 42348 6 wbs_dat_o[1]
port 197 nsew signal bidirectional
rlabel metal3 s 0 107388 800 107628 6 wbs_dat_o[20]
port 198 nsew signal bidirectional
rlabel metal3 s 0 164508 800 164748 6 wbs_dat_o[21]
port 199 nsew signal bidirectional
rlabel metal3 s 0 224348 800 224588 6 wbs_dat_o[22]
port 200 nsew signal bidirectional
rlabel metal3 s 0 79508 800 79748 6 wbs_dat_o[23]
port 201 nsew signal bidirectional
rlabel metal2 s 28970 0 29082 800 6 wbs_dat_o[24]
port 202 nsew signal bidirectional
rlabel metal2 s 10294 0 10406 800 6 wbs_dat_o[25]
port 203 nsew signal bidirectional
rlabel metal2 s 14802 239200 14914 240000 6 wbs_dat_o[26]
port 204 nsew signal bidirectional
rlabel metal3 s 0 221628 800 221868 6 wbs_dat_o[27]
port 205 nsew signal bidirectional
rlabel metal3 s 69200 8108 70000 8348 6 wbs_dat_o[28]
port 206 nsew signal bidirectional
rlabel metal2 s 36054 239200 36166 240000 6 wbs_dat_o[29]
port 207 nsew signal bidirectional
rlabel metal3 s 69200 118948 70000 119188 6 wbs_dat_o[2]
port 208 nsew signal bidirectional
rlabel metal3 s 0 118948 800 119188 6 wbs_dat_o[30]
port 209 nsew signal bidirectional
rlabel metal3 s 69200 195788 70000 196028 6 wbs_dat_o[31]
port 210 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 wbs_dat_o[3]
port 211 nsew signal bidirectional
rlabel metal2 s 53442 0 53554 800 6 wbs_dat_o[4]
port 212 nsew signal bidirectional
rlabel metal3 s 69200 16268 70000 16508 6 wbs_dat_o[5]
port 213 nsew signal bidirectional
rlabel metal3 s 69200 193068 70000 193308 6 wbs_dat_o[6]
port 214 nsew signal bidirectional
rlabel metal3 s 69200 18988 70000 19228 6 wbs_dat_o[7]
port 215 nsew signal bidirectional
rlabel metal2 s 25750 239200 25862 240000 6 wbs_dat_o[8]
port 216 nsew signal bidirectional
rlabel metal2 s 22530 239200 22642 240000 6 wbs_dat_o[9]
port 217 nsew signal bidirectional
rlabel metal3 s 0 150228 800 150468 6 wbs_sel_i[0]
port 218 nsew signal input
rlabel metal3 s 0 178788 800 179028 6 wbs_sel_i[1]
port 219 nsew signal input
rlabel metal3 s 69200 36668 70000 36908 6 wbs_sel_i[2]
port 220 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 wbs_sel_i[3]
port 221 nsew signal input
rlabel metal3 s 0 130508 800 130748 6 wbs_stb_i
port 222 nsew signal input
rlabel metal3 s 69200 158388 70000 158628 6 wbs_we_i
port 223 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 240000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 21054612
string GDS_FILE /home/runner/caravel_user_project/openlane/wrapped_etpu/runs/22_08_28_17_50/results/signoff/wrapped_etpu.magic.gds
string GDS_START 1011676
<< end >>

