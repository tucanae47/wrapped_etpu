magic
tech sky130A
magscale 1 2
timestamp 1654696751
<< obsli1 >>
rect 1104 2159 68816 69649
<< obsm1 >>
rect 14 2128 68816 69680
<< metal2 >>
rect 1278 71200 1390 72000
rect 3854 71200 3966 72000
rect 6430 71200 6542 72000
rect 9006 71200 9118 72000
rect 11582 71200 11694 72000
rect 14158 71200 14270 72000
rect 16734 71200 16846 72000
rect 19310 71200 19422 72000
rect 21886 71200 21998 72000
rect 24462 71200 24574 72000
rect 27038 71200 27150 72000
rect 29614 71200 29726 72000
rect 32190 71200 32302 72000
rect 34766 71200 34878 72000
rect 37342 71200 37454 72000
rect 39918 71200 40030 72000
rect 42494 71200 42606 72000
rect 45070 71200 45182 72000
rect 47646 71200 47758 72000
rect 50222 71200 50334 72000
rect 52798 71200 52910 72000
rect 55374 71200 55486 72000
rect 57950 71200 58062 72000
rect 60526 71200 60638 72000
rect 63102 71200 63214 72000
rect 65678 71200 65790 72000
rect 68254 71200 68366 72000
rect -10 0 102 800
rect 2566 0 2678 800
rect 5142 0 5254 800
rect 7718 0 7830 800
rect 10294 0 10406 800
rect 12870 0 12982 800
rect 15446 0 15558 800
rect 18022 0 18134 800
rect 20598 0 20710 800
rect 23174 0 23286 800
rect 25750 0 25862 800
rect 28326 0 28438 800
rect 30902 0 31014 800
rect 33478 0 33590 800
rect 36054 0 36166 800
rect 38630 0 38742 800
rect 41206 0 41318 800
rect 43782 0 43894 800
rect 46358 0 46470 800
rect 48934 0 49046 800
rect 51510 0 51622 800
rect 54086 0 54198 800
rect 56662 0 56774 800
rect 59238 0 59350 800
rect 61814 0 61926 800
rect 64390 0 64502 800
rect 66966 0 67078 800
rect 69542 0 69654 800
<< obsm2 >>
rect 20 71144 1222 71200
rect 1446 71144 3798 71200
rect 4022 71144 6374 71200
rect 6598 71144 8950 71200
rect 9174 71144 11526 71200
rect 11750 71144 14102 71200
rect 14326 71144 16678 71200
rect 16902 71144 19254 71200
rect 19478 71144 21830 71200
rect 22054 71144 24406 71200
rect 24630 71144 26982 71200
rect 27206 71144 29558 71200
rect 29782 71144 32134 71200
rect 32358 71144 34710 71200
rect 34934 71144 37286 71200
rect 37510 71144 39862 71200
rect 40086 71144 42438 71200
rect 42662 71144 45014 71200
rect 45238 71144 47590 71200
rect 47814 71144 50166 71200
rect 50390 71144 52742 71200
rect 52966 71144 55318 71200
rect 55542 71144 57894 71200
rect 58118 71144 60470 71200
rect 60694 71144 63046 71200
rect 63270 71144 65622 71200
rect 65846 71144 68198 71200
rect 20 856 68336 71144
rect 158 734 2510 856
rect 2734 734 5086 856
rect 5310 734 7662 856
rect 7886 734 10238 856
rect 10462 734 12814 856
rect 13038 734 15390 856
rect 15614 734 17966 856
rect 18190 734 20542 856
rect 20766 734 23118 856
rect 23342 734 25694 856
rect 25918 734 28270 856
rect 28494 734 30846 856
rect 31070 734 33422 856
rect 33646 734 35998 856
rect 36222 734 38574 856
rect 38798 734 41150 856
rect 41374 734 43726 856
rect 43950 734 46302 856
rect 46526 734 48878 856
rect 49102 734 51454 856
rect 51678 734 54030 856
rect 54254 734 56606 856
rect 56830 734 59182 856
rect 59406 734 61758 856
rect 61982 734 64334 856
rect 64558 734 66910 856
rect 67134 734 68336 856
<< metal3 >>
rect 0 70668 800 70908
rect 69200 69988 70000 70228
rect 0 67948 800 68188
rect 69200 67268 70000 67508
rect 0 65228 800 65468
rect 69200 64548 70000 64788
rect 0 62508 800 62748
rect 69200 61828 70000 62068
rect 0 59788 800 60028
rect 69200 59108 70000 59348
rect 0 57068 800 57308
rect 69200 56388 70000 56628
rect 0 54348 800 54588
rect 69200 53668 70000 53908
rect 0 51628 800 51868
rect 69200 50948 70000 51188
rect 0 48908 800 49148
rect 69200 48228 70000 48468
rect 0 46188 800 46428
rect 69200 45508 70000 45748
rect 0 43468 800 43708
rect 69200 42788 70000 43028
rect 0 40748 800 40988
rect 69200 40068 70000 40308
rect 0 38028 800 38268
rect 69200 37348 70000 37588
rect 0 35308 800 35548
rect 69200 34628 70000 34868
rect 0 32588 800 32828
rect 69200 31908 70000 32148
rect 0 29868 800 30108
rect 69200 29188 70000 29428
rect 0 27148 800 27388
rect 69200 26468 70000 26708
rect 0 24428 800 24668
rect 69200 23748 70000 23988
rect 0 21708 800 21948
rect 69200 21028 70000 21268
rect 0 18988 800 19228
rect 69200 18308 70000 18548
rect 0 16268 800 16508
rect 69200 15588 70000 15828
rect 0 13548 800 13788
rect 69200 12868 70000 13108
rect 0 10828 800 11068
rect 69200 10148 70000 10388
rect 0 8108 800 8348
rect 69200 7428 70000 7668
rect 0 5388 800 5628
rect 69200 4708 70000 4948
rect 0 2668 800 2908
rect 69200 1988 70000 2228
<< obsm3 >>
rect 880 70588 69200 70821
rect 800 70308 69200 70588
rect 800 69908 69120 70308
rect 800 68268 69200 69908
rect 880 67868 69200 68268
rect 800 67588 69200 67868
rect 800 67188 69120 67588
rect 800 65548 69200 67188
rect 880 65148 69200 65548
rect 800 64868 69200 65148
rect 800 64468 69120 64868
rect 800 62828 69200 64468
rect 880 62428 69200 62828
rect 800 62148 69200 62428
rect 800 61748 69120 62148
rect 800 60108 69200 61748
rect 880 59708 69200 60108
rect 800 59428 69200 59708
rect 800 59028 69120 59428
rect 800 57388 69200 59028
rect 880 56988 69200 57388
rect 800 56708 69200 56988
rect 800 56308 69120 56708
rect 800 54668 69200 56308
rect 880 54268 69200 54668
rect 800 53988 69200 54268
rect 800 53588 69120 53988
rect 800 51948 69200 53588
rect 880 51548 69200 51948
rect 800 51268 69200 51548
rect 800 50868 69120 51268
rect 800 49228 69200 50868
rect 880 48828 69200 49228
rect 800 48548 69200 48828
rect 800 48148 69120 48548
rect 800 46508 69200 48148
rect 880 46108 69200 46508
rect 800 45828 69200 46108
rect 800 45428 69120 45828
rect 800 43788 69200 45428
rect 880 43388 69200 43788
rect 800 43108 69200 43388
rect 800 42708 69120 43108
rect 800 41068 69200 42708
rect 880 40668 69200 41068
rect 800 40388 69200 40668
rect 800 39988 69120 40388
rect 800 38348 69200 39988
rect 880 37948 69200 38348
rect 800 37668 69200 37948
rect 800 37268 69120 37668
rect 800 35628 69200 37268
rect 880 35228 69200 35628
rect 800 34948 69200 35228
rect 800 34548 69120 34948
rect 800 32908 69200 34548
rect 880 32508 69200 32908
rect 800 32228 69200 32508
rect 800 31828 69120 32228
rect 800 30188 69200 31828
rect 880 29788 69200 30188
rect 800 29508 69200 29788
rect 800 29108 69120 29508
rect 800 27468 69200 29108
rect 880 27068 69200 27468
rect 800 26788 69200 27068
rect 800 26388 69120 26788
rect 800 24748 69200 26388
rect 880 24348 69200 24748
rect 800 24068 69200 24348
rect 800 23668 69120 24068
rect 800 22028 69200 23668
rect 880 21628 69200 22028
rect 800 21348 69200 21628
rect 800 20948 69120 21348
rect 800 19308 69200 20948
rect 880 18908 69200 19308
rect 800 18628 69200 18908
rect 800 18228 69120 18628
rect 800 16588 69200 18228
rect 880 16188 69200 16588
rect 800 15908 69200 16188
rect 800 15508 69120 15908
rect 800 13868 69200 15508
rect 880 13468 69200 13868
rect 800 13188 69200 13468
rect 800 12788 69120 13188
rect 800 11148 69200 12788
rect 880 10748 69200 11148
rect 800 10468 69200 10748
rect 800 10068 69120 10468
rect 800 8428 69200 10068
rect 880 8028 69200 8428
rect 800 7748 69200 8028
rect 800 7348 69120 7748
rect 800 5708 69200 7348
rect 880 5308 69200 5708
rect 800 5028 69200 5308
rect 800 4628 69120 5028
rect 800 2988 69200 4628
rect 880 2588 69200 2988
rect 800 2308 69200 2588
rect 800 2143 69120 2308
<< metal4 >>
rect 4208 2128 4528 69680
rect 19568 2128 19888 69680
rect 34928 2128 35248 69680
rect 50288 2128 50608 69680
rect 65648 2128 65968 69680
<< labels >>
rlabel metal3 s 0 70668 800 70908 6 active
port 1 nsew signal input
rlabel metal4 s 4208 2128 4528 69680 6 vccd1
port 2 nsew power input
rlabel metal4 s 34928 2128 35248 69680 6 vccd1
port 2 nsew power input
rlabel metal4 s 65648 2128 65968 69680 6 vccd1
port 2 nsew power input
rlabel metal4 s 19568 2128 19888 69680 6 vssd1
port 3 nsew ground input
rlabel metal4 s 50288 2128 50608 69680 6 vssd1
port 3 nsew ground input
rlabel metal3 s 69200 69988 70000 70228 6 wb_clk_i
port 4 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 wb_rst_i
port 5 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 wbs_ack_o
port 6 nsew signal bidirectional
rlabel metal3 s 0 40748 800 40988 6 wbs_adr_i[0]
port 7 nsew signal input
rlabel metal2 s 42494 71200 42606 72000 6 wbs_adr_i[10]
port 8 nsew signal input
rlabel metal2 s 65678 71200 65790 72000 6 wbs_adr_i[11]
port 9 nsew signal input
rlabel metal2 s 50222 71200 50334 72000 6 wbs_adr_i[12]
port 10 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 wbs_adr_i[13]
port 11 nsew signal input
rlabel metal2 s 34766 71200 34878 72000 6 wbs_adr_i[14]
port 12 nsew signal input
rlabel metal2 s 64390 0 64502 800 6 wbs_adr_i[15]
port 13 nsew signal input
rlabel metal3 s 69200 40068 70000 40308 6 wbs_adr_i[16]
port 14 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 wbs_adr_i[17]
port 15 nsew signal input
rlabel metal3 s 0 54348 800 54588 6 wbs_adr_i[18]
port 16 nsew signal input
rlabel metal2 s 47646 71200 47758 72000 6 wbs_adr_i[19]
port 17 nsew signal input
rlabel metal2 s 61814 0 61926 800 6 wbs_adr_i[1]
port 18 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 wbs_adr_i[20]
port 19 nsew signal input
rlabel metal3 s 69200 61828 70000 62068 6 wbs_adr_i[21]
port 20 nsew signal input
rlabel metal3 s 0 59788 800 60028 6 wbs_adr_i[22]
port 21 nsew signal input
rlabel metal3 s 69200 23748 70000 23988 6 wbs_adr_i[23]
port 22 nsew signal input
rlabel metal3 s 69200 59108 70000 59348 6 wbs_adr_i[24]
port 23 nsew signal input
rlabel metal2 s 57950 71200 58062 72000 6 wbs_adr_i[25]
port 24 nsew signal input
rlabel metal3 s 69200 15588 70000 15828 6 wbs_adr_i[26]
port 25 nsew signal input
rlabel metal3 s 69200 67268 70000 67508 6 wbs_adr_i[27]
port 26 nsew signal input
rlabel metal3 s 0 13548 800 13788 6 wbs_adr_i[28]
port 27 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 wbs_adr_i[29]
port 28 nsew signal input
rlabel metal3 s 69200 12868 70000 13108 6 wbs_adr_i[2]
port 29 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 wbs_adr_i[30]
port 30 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 wbs_adr_i[31]
port 31 nsew signal input
rlabel metal2 s 19310 71200 19422 72000 6 wbs_adr_i[3]
port 32 nsew signal input
rlabel metal2 s 37342 71200 37454 72000 6 wbs_adr_i[4]
port 33 nsew signal input
rlabel metal2 s 63102 71200 63214 72000 6 wbs_adr_i[5]
port 34 nsew signal input
rlabel metal2 s 7718 0 7830 800 6 wbs_adr_i[6]
port 35 nsew signal input
rlabel metal3 s 69200 53668 70000 53908 6 wbs_adr_i[7]
port 36 nsew signal input
rlabel metal3 s 0 46188 800 46428 6 wbs_adr_i[8]
port 37 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 wbs_adr_i[9]
port 38 nsew signal input
rlabel metal3 s 69200 4708 70000 4948 6 wbs_cyc_i
port 39 nsew signal input
rlabel metal2 s 54086 0 54198 800 6 wbs_dat_i[0]
port 40 nsew signal input
rlabel metal3 s 69200 31908 70000 32148 6 wbs_dat_i[10]
port 41 nsew signal input
rlabel metal3 s 69200 26468 70000 26708 6 wbs_dat_i[11]
port 42 nsew signal input
rlabel metal2 s 21886 71200 21998 72000 6 wbs_dat_i[12]
port 43 nsew signal input
rlabel metal2 s 24462 71200 24574 72000 6 wbs_dat_i[13]
port 44 nsew signal input
rlabel metal3 s 69200 56388 70000 56628 6 wbs_dat_i[14]
port 45 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 wbs_dat_i[15]
port 46 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 wbs_dat_i[16]
port 47 nsew signal input
rlabel metal3 s 69200 10148 70000 10388 6 wbs_dat_i[17]
port 48 nsew signal input
rlabel metal3 s 69200 1988 70000 2228 6 wbs_dat_i[18]
port 49 nsew signal input
rlabel metal3 s 69200 37348 70000 37588 6 wbs_dat_i[19]
port 50 nsew signal input
rlabel metal3 s 0 51628 800 51868 6 wbs_dat_i[1]
port 51 nsew signal input
rlabel metal2 s 59238 0 59350 800 6 wbs_dat_i[20]
port 52 nsew signal input
rlabel metal2 s 27038 71200 27150 72000 6 wbs_dat_i[21]
port 53 nsew signal input
rlabel metal3 s 69200 64548 70000 64788 6 wbs_dat_i[22]
port 54 nsew signal input
rlabel metal2 s 69542 0 69654 800 6 wbs_dat_i[23]
port 55 nsew signal input
rlabel metal2 s 32190 71200 32302 72000 6 wbs_dat_i[24]
port 56 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 wbs_dat_i[25]
port 57 nsew signal input
rlabel metal3 s 69200 18308 70000 18548 6 wbs_dat_i[26]
port 58 nsew signal input
rlabel metal3 s 69200 45508 70000 45748 6 wbs_dat_i[27]
port 59 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 wbs_dat_i[28]
port 60 nsew signal input
rlabel metal2 s 39918 71200 40030 72000 6 wbs_dat_i[29]
port 61 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 wbs_dat_i[2]
port 62 nsew signal input
rlabel metal2 s 16734 71200 16846 72000 6 wbs_dat_i[30]
port 63 nsew signal input
rlabel metal3 s 0 65228 800 65468 6 wbs_dat_i[31]
port 64 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 wbs_dat_i[3]
port 65 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 wbs_dat_i[4]
port 66 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 wbs_dat_i[5]
port 67 nsew signal input
rlabel metal2 s 66966 0 67078 800 6 wbs_dat_i[6]
port 68 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 wbs_dat_i[7]
port 69 nsew signal input
rlabel metal3 s 69200 21028 70000 21268 6 wbs_dat_i[8]
port 70 nsew signal input
rlabel metal2 s 51510 0 51622 800 6 wbs_dat_i[9]
port 71 nsew signal input
rlabel metal3 s 0 57068 800 57308 6 wbs_dat_o[0]
port 72 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 wbs_dat_o[10]
port 73 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 wbs_dat_o[11]
port 74 nsew signal bidirectional
rlabel metal3 s 69200 29188 70000 29428 6 wbs_dat_o[12]
port 75 nsew signal bidirectional
rlabel metal3 s 69200 48228 70000 48468 6 wbs_dat_o[13]
port 76 nsew signal bidirectional
rlabel metal2 s 56662 0 56774 800 6 wbs_dat_o[14]
port 77 nsew signal bidirectional
rlabel metal3 s 69200 50948 70000 51188 6 wbs_dat_o[15]
port 78 nsew signal bidirectional
rlabel metal2 s 6430 71200 6542 72000 6 wbs_dat_o[16]
port 79 nsew signal bidirectional
rlabel metal2 s 9006 71200 9118 72000 6 wbs_dat_o[17]
port 80 nsew signal bidirectional
rlabel metal2 s 36054 0 36166 800 6 wbs_dat_o[18]
port 81 nsew signal bidirectional
rlabel metal2 s -10 0 102 800 6 wbs_dat_o[19]
port 82 nsew signal bidirectional
rlabel metal2 s 43782 0 43894 800 6 wbs_dat_o[1]
port 83 nsew signal bidirectional
rlabel metal2 s 11582 71200 11694 72000 6 wbs_dat_o[20]
port 84 nsew signal bidirectional
rlabel metal2 s 29614 71200 29726 72000 6 wbs_dat_o[21]
port 85 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 wbs_dat_o[22]
port 86 nsew signal bidirectional
rlabel metal3 s 0 67948 800 68188 6 wbs_dat_o[23]
port 87 nsew signal bidirectional
rlabel metal2 s 10294 0 10406 800 6 wbs_dat_o[24]
port 88 nsew signal bidirectional
rlabel metal2 s 2566 0 2678 800 6 wbs_dat_o[25]
port 89 nsew signal bidirectional
rlabel metal2 s 60526 71200 60638 72000 6 wbs_dat_o[26]
port 90 nsew signal bidirectional
rlabel metal2 s 45070 71200 45182 72000 6 wbs_dat_o[27]
port 91 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 wbs_dat_o[28]
port 92 nsew signal bidirectional
rlabel metal2 s 68254 71200 68366 72000 6 wbs_dat_o[29]
port 93 nsew signal bidirectional
rlabel metal3 s 69200 7428 70000 7668 6 wbs_dat_o[2]
port 94 nsew signal bidirectional
rlabel metal2 s 1278 71200 1390 72000 6 wbs_dat_o[30]
port 95 nsew signal bidirectional
rlabel metal3 s 0 27148 800 27388 6 wbs_dat_o[31]
port 96 nsew signal bidirectional
rlabel metal2 s 12870 0 12982 800 6 wbs_dat_o[3]
port 97 nsew signal bidirectional
rlabel metal2 s 23174 0 23286 800 6 wbs_dat_o[4]
port 98 nsew signal bidirectional
rlabel metal3 s 0 24428 800 24668 6 wbs_dat_o[5]
port 99 nsew signal bidirectional
rlabel metal3 s 69200 42788 70000 43028 6 wbs_dat_o[6]
port 100 nsew signal bidirectional
rlabel metal2 s 38630 0 38742 800 6 wbs_dat_o[7]
port 101 nsew signal bidirectional
rlabel metal2 s 55374 71200 55486 72000 6 wbs_dat_o[8]
port 102 nsew signal bidirectional
rlabel metal2 s 52798 71200 52910 72000 6 wbs_dat_o[9]
port 103 nsew signal bidirectional
rlabel metal2 s 3854 71200 3966 72000 6 wbs_sel_i[0]
port 104 nsew signal input
rlabel metal2 s 14158 71200 14270 72000 6 wbs_sel_i[1]
port 105 nsew signal input
rlabel metal2 s 48934 0 49046 800 6 wbs_sel_i[2]
port 106 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 wbs_sel_i[3]
port 107 nsew signal input
rlabel metal3 s 0 62508 800 62748 6 wbs_stb_i
port 108 nsew signal input
rlabel metal3 s 69200 34628 70000 34868 6 wbs_we_i
port 109 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 72000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1612790
string GDS_FILE /home/tuc/MPW5/caravel_user_project/openlane/wrapped_etpu/runs/wrapped_etpu/results/finishing/wrapped_etpu.magic.gds
string GDS_START 138124
<< end >>

