magic
tech sky130B
magscale 1 2
timestamp 1661706560
<< obsli1 >>
rect 1104 2159 178848 177361
<< obsm1 >>
rect 14 1300 178848 177392
<< metal2 >>
rect 634 179200 746 180000
rect 3854 179200 3966 180000
rect 7074 179200 7186 180000
rect 10294 179200 10406 180000
rect 13514 179200 13626 180000
rect 16090 179200 16202 180000
rect 19310 179200 19422 180000
rect 22530 179200 22642 180000
rect 25750 179200 25862 180000
rect 28970 179200 29082 180000
rect 32190 179200 32302 180000
rect 35410 179200 35522 180000
rect 38630 179200 38742 180000
rect 41850 179200 41962 180000
rect 45070 179200 45182 180000
rect 48290 179200 48402 180000
rect 51510 179200 51622 180000
rect 54730 179200 54842 180000
rect 57950 179200 58062 180000
rect 61170 179200 61282 180000
rect 63746 179200 63858 180000
rect 66966 179200 67078 180000
rect 70186 179200 70298 180000
rect 73406 179200 73518 180000
rect 76626 179200 76738 180000
rect 79846 179200 79958 180000
rect 83066 179200 83178 180000
rect 86286 179200 86398 180000
rect 89506 179200 89618 180000
rect 92726 179200 92838 180000
rect 95946 179200 96058 180000
rect 99166 179200 99278 180000
rect 102386 179200 102498 180000
rect 105606 179200 105718 180000
rect 108826 179200 108938 180000
rect 111402 179200 111514 180000
rect 114622 179200 114734 180000
rect 117842 179200 117954 180000
rect 121062 179200 121174 180000
rect 124282 179200 124394 180000
rect 127502 179200 127614 180000
rect 130722 179200 130834 180000
rect 133942 179200 134054 180000
rect 137162 179200 137274 180000
rect 140382 179200 140494 180000
rect 143602 179200 143714 180000
rect 146822 179200 146934 180000
rect 150042 179200 150154 180000
rect 153262 179200 153374 180000
rect 156482 179200 156594 180000
rect 159058 179200 159170 180000
rect 162278 179200 162390 180000
rect 165498 179200 165610 180000
rect 168718 179200 168830 180000
rect 171938 179200 172050 180000
rect 175158 179200 175270 180000
rect 178378 179200 178490 180000
rect -10 0 102 800
rect 2566 0 2678 800
rect 5786 0 5898 800
rect 9006 0 9118 800
rect 12226 0 12338 800
rect 15446 0 15558 800
rect 18666 0 18778 800
rect 21886 0 21998 800
rect 25106 0 25218 800
rect 28326 0 28438 800
rect 31546 0 31658 800
rect 34766 0 34878 800
rect 37986 0 38098 800
rect 41206 0 41318 800
rect 44426 0 44538 800
rect 47002 0 47114 800
rect 50222 0 50334 800
rect 53442 0 53554 800
rect 56662 0 56774 800
rect 59882 0 59994 800
rect 63102 0 63214 800
rect 66322 0 66434 800
rect 69542 0 69654 800
rect 72762 0 72874 800
rect 75982 0 76094 800
rect 79202 0 79314 800
rect 82422 0 82534 800
rect 85642 0 85754 800
rect 88862 0 88974 800
rect 92082 0 92194 800
rect 94658 0 94770 800
rect 97878 0 97990 800
rect 101098 0 101210 800
rect 104318 0 104430 800
rect 107538 0 107650 800
rect 110758 0 110870 800
rect 113978 0 114090 800
rect 117198 0 117310 800
rect 120418 0 120530 800
rect 123638 0 123750 800
rect 126858 0 126970 800
rect 130078 0 130190 800
rect 133298 0 133410 800
rect 136518 0 136630 800
rect 139738 0 139850 800
rect 142314 0 142426 800
rect 145534 0 145646 800
rect 148754 0 148866 800
rect 151974 0 152086 800
rect 155194 0 155306 800
rect 158414 0 158526 800
rect 161634 0 161746 800
rect 164854 0 164966 800
rect 168074 0 168186 800
rect 171294 0 171406 800
rect 174514 0 174626 800
rect 177734 0 177846 800
<< obsm2 >>
rect 20 179144 578 179466
rect 802 179144 3798 179466
rect 4022 179144 7018 179466
rect 7242 179144 10238 179466
rect 10462 179144 13458 179466
rect 13682 179144 16034 179466
rect 16258 179144 19254 179466
rect 19478 179144 22474 179466
rect 22698 179144 25694 179466
rect 25918 179144 28914 179466
rect 29138 179144 32134 179466
rect 32358 179144 35354 179466
rect 35578 179144 38574 179466
rect 38798 179144 41794 179466
rect 42018 179144 45014 179466
rect 45238 179144 48234 179466
rect 48458 179144 51454 179466
rect 51678 179144 54674 179466
rect 54898 179144 57894 179466
rect 58118 179144 61114 179466
rect 61338 179144 63690 179466
rect 63914 179144 66910 179466
rect 67134 179144 70130 179466
rect 70354 179144 73350 179466
rect 73574 179144 76570 179466
rect 76794 179144 79790 179466
rect 80014 179144 83010 179466
rect 83234 179144 86230 179466
rect 86454 179144 89450 179466
rect 89674 179144 92670 179466
rect 92894 179144 95890 179466
rect 96114 179144 99110 179466
rect 99334 179144 102330 179466
rect 102554 179144 105550 179466
rect 105774 179144 108770 179466
rect 108994 179144 111346 179466
rect 111570 179144 114566 179466
rect 114790 179144 117786 179466
rect 118010 179144 121006 179466
rect 121230 179144 124226 179466
rect 124450 179144 127446 179466
rect 127670 179144 130666 179466
rect 130890 179144 133886 179466
rect 134110 179144 137106 179466
rect 137330 179144 140326 179466
rect 140550 179144 143546 179466
rect 143770 179144 146766 179466
rect 146990 179144 149986 179466
rect 150210 179144 153206 179466
rect 153430 179144 156426 179466
rect 156650 179144 159002 179466
rect 159226 179144 162222 179466
rect 162446 179144 165442 179466
rect 165666 179144 168662 179466
rect 168886 179144 171882 179466
rect 172106 179144 175102 179466
rect 175326 179144 178322 179466
rect 20 856 178460 179144
rect 158 711 2510 856
rect 2734 711 5730 856
rect 5954 711 8950 856
rect 9174 711 12170 856
rect 12394 711 15390 856
rect 15614 711 18610 856
rect 18834 711 21830 856
rect 22054 711 25050 856
rect 25274 711 28270 856
rect 28494 711 31490 856
rect 31714 711 34710 856
rect 34934 711 37930 856
rect 38154 711 41150 856
rect 41374 711 44370 856
rect 44594 711 46946 856
rect 47170 711 50166 856
rect 50390 711 53386 856
rect 53610 711 56606 856
rect 56830 711 59826 856
rect 60050 711 63046 856
rect 63270 711 66266 856
rect 66490 711 69486 856
rect 69710 711 72706 856
rect 72930 711 75926 856
rect 76150 711 79146 856
rect 79370 711 82366 856
rect 82590 711 85586 856
rect 85810 711 88806 856
rect 89030 711 92026 856
rect 92250 711 94602 856
rect 94826 711 97822 856
rect 98046 711 101042 856
rect 101266 711 104262 856
rect 104486 711 107482 856
rect 107706 711 110702 856
rect 110926 711 113922 856
rect 114146 711 117142 856
rect 117366 711 120362 856
rect 120586 711 123582 856
rect 123806 711 126802 856
rect 127026 711 130022 856
rect 130246 711 133242 856
rect 133466 711 136462 856
rect 136686 711 139682 856
rect 139906 711 142258 856
rect 142482 711 145478 856
rect 145702 711 148698 856
rect 148922 711 151918 856
rect 152142 711 155138 856
rect 155362 711 158358 856
rect 158582 711 161578 856
rect 161802 711 164798 856
rect 165022 711 168018 856
rect 168242 711 171238 856
rect 171462 711 174458 856
rect 174682 711 177678 856
rect 177902 711 178460 856
<< metal3 >>
rect 179200 178108 180000 178348
rect 0 177428 800 177668
rect 179200 174708 180000 174948
rect 0 174028 800 174268
rect 179200 171308 180000 171548
rect 0 170628 800 170868
rect 179200 167908 180000 168148
rect 0 167228 800 167468
rect 179200 164508 180000 164748
rect 0 163828 800 164068
rect 179200 161108 180000 161348
rect 0 160428 800 160668
rect 179200 157708 180000 157948
rect 0 157028 800 157268
rect 179200 154988 180000 155228
rect 0 153628 800 153868
rect 179200 151588 180000 151828
rect 0 150228 800 150468
rect 179200 148188 180000 148428
rect 0 147508 800 147748
rect 179200 144788 180000 145028
rect 0 144108 800 144348
rect 179200 141388 180000 141628
rect 0 140708 800 140948
rect 179200 137988 180000 138228
rect 0 137308 800 137548
rect 179200 134588 180000 134828
rect 0 133908 800 134148
rect 179200 131188 180000 131428
rect 0 130508 800 130748
rect 179200 127788 180000 128028
rect 0 127108 800 127348
rect 179200 124388 180000 124628
rect 0 123708 800 123948
rect 179200 120988 180000 121228
rect 0 120308 800 120548
rect 179200 117588 180000 117828
rect 0 116908 800 117148
rect 179200 114188 180000 114428
rect 0 113508 800 113748
rect 179200 110788 180000 111028
rect 0 110108 800 110348
rect 179200 107388 180000 107628
rect 0 106708 800 106948
rect 179200 104668 180000 104908
rect 0 103308 800 103548
rect 179200 101268 180000 101508
rect 0 99908 800 100148
rect 179200 97868 180000 98108
rect 0 97188 800 97428
rect 179200 94468 180000 94708
rect 0 93788 800 94028
rect 179200 91068 180000 91308
rect 0 90388 800 90628
rect 179200 87668 180000 87908
rect 0 86988 800 87228
rect 179200 84268 180000 84508
rect 0 83588 800 83828
rect 179200 80868 180000 81108
rect 0 80188 800 80428
rect 179200 77468 180000 77708
rect 0 76788 800 77028
rect 179200 74068 180000 74308
rect 0 73388 800 73628
rect 179200 70668 180000 70908
rect 0 69988 800 70228
rect 179200 67268 180000 67508
rect 0 66588 800 66828
rect 179200 63868 180000 64108
rect 0 63188 800 63428
rect 179200 60468 180000 60708
rect 0 59788 800 60028
rect 179200 57068 180000 57308
rect 0 56388 800 56628
rect 179200 54348 180000 54588
rect 0 52988 800 53228
rect 179200 50948 180000 51188
rect 0 49588 800 49828
rect 179200 47548 180000 47788
rect 0 46868 800 47108
rect 179200 44148 180000 44388
rect 0 43468 800 43708
rect 179200 40748 180000 40988
rect 0 40068 800 40308
rect 179200 37348 180000 37588
rect 0 36668 800 36908
rect 179200 33948 180000 34188
rect 0 33268 800 33508
rect 179200 30548 180000 30788
rect 0 29868 800 30108
rect 179200 27148 180000 27388
rect 0 26468 800 26708
rect 179200 23748 180000 23988
rect 0 23068 800 23308
rect 179200 20348 180000 20588
rect 0 19668 800 19908
rect 179200 16948 180000 17188
rect 0 16268 800 16508
rect 179200 13548 180000 13788
rect 0 12868 800 13108
rect 179200 10148 180000 10388
rect 0 9468 800 9708
rect 179200 6748 180000 6988
rect 0 6068 800 6308
rect 179200 4028 180000 4268
rect 0 2668 800 2908
rect 179200 628 180000 868
<< obsm3 >>
rect 800 178028 179120 178261
rect 800 177748 179200 178028
rect 880 177348 179200 177748
rect 800 175028 179200 177348
rect 800 174628 179120 175028
rect 800 174348 179200 174628
rect 880 173948 179200 174348
rect 800 171628 179200 173948
rect 800 171228 179120 171628
rect 800 170948 179200 171228
rect 880 170548 179200 170948
rect 800 168228 179200 170548
rect 800 167828 179120 168228
rect 800 167548 179200 167828
rect 880 167148 179200 167548
rect 800 164828 179200 167148
rect 800 164428 179120 164828
rect 800 164148 179200 164428
rect 880 163748 179200 164148
rect 800 161428 179200 163748
rect 800 161028 179120 161428
rect 800 160748 179200 161028
rect 880 160348 179200 160748
rect 800 158028 179200 160348
rect 800 157628 179120 158028
rect 800 157348 179200 157628
rect 880 156948 179200 157348
rect 800 155308 179200 156948
rect 800 154908 179120 155308
rect 800 153948 179200 154908
rect 880 153548 179200 153948
rect 800 151908 179200 153548
rect 800 151508 179120 151908
rect 800 150548 179200 151508
rect 880 150148 179200 150548
rect 800 148508 179200 150148
rect 800 148108 179120 148508
rect 800 147828 179200 148108
rect 880 147428 179200 147828
rect 800 145108 179200 147428
rect 800 144708 179120 145108
rect 800 144428 179200 144708
rect 880 144028 179200 144428
rect 800 141708 179200 144028
rect 800 141308 179120 141708
rect 800 141028 179200 141308
rect 880 140628 179200 141028
rect 800 138308 179200 140628
rect 800 137908 179120 138308
rect 800 137628 179200 137908
rect 880 137228 179200 137628
rect 800 134908 179200 137228
rect 800 134508 179120 134908
rect 800 134228 179200 134508
rect 880 133828 179200 134228
rect 800 131508 179200 133828
rect 800 131108 179120 131508
rect 800 130828 179200 131108
rect 880 130428 179200 130828
rect 800 128108 179200 130428
rect 800 127708 179120 128108
rect 800 127428 179200 127708
rect 880 127028 179200 127428
rect 800 124708 179200 127028
rect 800 124308 179120 124708
rect 800 124028 179200 124308
rect 880 123628 179200 124028
rect 800 121308 179200 123628
rect 800 120908 179120 121308
rect 800 120628 179200 120908
rect 880 120228 179200 120628
rect 800 117908 179200 120228
rect 800 117508 179120 117908
rect 800 117228 179200 117508
rect 880 116828 179200 117228
rect 800 114508 179200 116828
rect 800 114108 179120 114508
rect 800 113828 179200 114108
rect 880 113428 179200 113828
rect 800 111108 179200 113428
rect 800 110708 179120 111108
rect 800 110428 179200 110708
rect 880 110028 179200 110428
rect 800 107708 179200 110028
rect 800 107308 179120 107708
rect 800 107028 179200 107308
rect 880 106628 179200 107028
rect 800 104988 179200 106628
rect 800 104588 179120 104988
rect 800 103628 179200 104588
rect 880 103228 179200 103628
rect 800 101588 179200 103228
rect 800 101188 179120 101588
rect 800 100228 179200 101188
rect 880 99828 179200 100228
rect 800 98188 179200 99828
rect 800 97788 179120 98188
rect 800 97508 179200 97788
rect 880 97108 179200 97508
rect 800 94788 179200 97108
rect 800 94388 179120 94788
rect 800 94108 179200 94388
rect 880 93708 179200 94108
rect 800 91388 179200 93708
rect 800 90988 179120 91388
rect 800 90708 179200 90988
rect 880 90308 179200 90708
rect 800 87988 179200 90308
rect 800 87588 179120 87988
rect 800 87308 179200 87588
rect 880 86908 179200 87308
rect 800 84588 179200 86908
rect 800 84188 179120 84588
rect 800 83908 179200 84188
rect 880 83508 179200 83908
rect 800 81188 179200 83508
rect 800 80788 179120 81188
rect 800 80508 179200 80788
rect 880 80108 179200 80508
rect 800 77788 179200 80108
rect 800 77388 179120 77788
rect 800 77108 179200 77388
rect 880 76708 179200 77108
rect 800 74388 179200 76708
rect 800 73988 179120 74388
rect 800 73708 179200 73988
rect 880 73308 179200 73708
rect 800 70988 179200 73308
rect 800 70588 179120 70988
rect 800 70308 179200 70588
rect 880 69908 179200 70308
rect 800 67588 179200 69908
rect 800 67188 179120 67588
rect 800 66908 179200 67188
rect 880 66508 179200 66908
rect 800 64188 179200 66508
rect 800 63788 179120 64188
rect 800 63508 179200 63788
rect 880 63108 179200 63508
rect 800 60788 179200 63108
rect 800 60388 179120 60788
rect 800 60108 179200 60388
rect 880 59708 179200 60108
rect 800 57388 179200 59708
rect 800 56988 179120 57388
rect 800 56708 179200 56988
rect 880 56308 179200 56708
rect 800 54668 179200 56308
rect 800 54268 179120 54668
rect 800 53308 179200 54268
rect 880 52908 179200 53308
rect 800 51268 179200 52908
rect 800 50868 179120 51268
rect 800 49908 179200 50868
rect 880 49508 179200 49908
rect 800 47868 179200 49508
rect 800 47468 179120 47868
rect 800 47188 179200 47468
rect 880 46788 179200 47188
rect 800 44468 179200 46788
rect 800 44068 179120 44468
rect 800 43788 179200 44068
rect 880 43388 179200 43788
rect 800 41068 179200 43388
rect 800 40668 179120 41068
rect 800 40388 179200 40668
rect 880 39988 179200 40388
rect 800 37668 179200 39988
rect 800 37268 179120 37668
rect 800 36988 179200 37268
rect 880 36588 179200 36988
rect 800 34268 179200 36588
rect 800 33868 179120 34268
rect 800 33588 179200 33868
rect 880 33188 179200 33588
rect 800 30868 179200 33188
rect 800 30468 179120 30868
rect 800 30188 179200 30468
rect 880 29788 179200 30188
rect 800 27468 179200 29788
rect 800 27068 179120 27468
rect 800 26788 179200 27068
rect 880 26388 179200 26788
rect 800 24068 179200 26388
rect 800 23668 179120 24068
rect 800 23388 179200 23668
rect 880 22988 179200 23388
rect 800 20668 179200 22988
rect 800 20268 179120 20668
rect 800 19988 179200 20268
rect 880 19588 179200 19988
rect 800 17268 179200 19588
rect 800 16868 179120 17268
rect 800 16588 179200 16868
rect 880 16188 179200 16588
rect 800 13868 179200 16188
rect 800 13468 179120 13868
rect 800 13188 179200 13468
rect 880 12788 179200 13188
rect 800 10468 179200 12788
rect 800 10068 179120 10468
rect 800 9788 179200 10068
rect 880 9388 179200 9788
rect 800 7068 179200 9388
rect 800 6668 179120 7068
rect 800 6388 179200 6668
rect 880 5988 179200 6388
rect 800 4348 179200 5988
rect 800 3948 179120 4348
rect 800 2988 179200 3948
rect 880 2588 179200 2988
rect 800 948 179200 2588
rect 800 715 179120 948
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
<< obsm4 >>
rect 50843 2347 65568 150517
rect 66048 2347 80928 150517
rect 81408 2347 96288 150517
rect 96768 2347 111648 150517
rect 112128 2347 127008 150517
rect 127488 2347 142368 150517
rect 142848 2347 153397 150517
<< labels >>
rlabel metal2 s 634 179200 746 180000 6 active
port 1 nsew signal input
rlabel metal3 s 179200 54348 180000 54588 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 133298 0 133410 800 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 139738 0 139850 800 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 io_in[12]
port 5 nsew signal input
rlabel metal3 s 179200 27148 180000 27388 6 io_in[13]
port 6 nsew signal input
rlabel metal3 s 179200 20348 180000 20588 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 66322 0 66434 800 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 179200 91068 180000 91308 6 io_in[17]
port 10 nsew signal input
rlabel metal3 s 179200 67268 180000 67508 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 145534 0 145646 800 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 57950 179200 58062 180000 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 179200 4028 180000 4268 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 179200 131188 180000 131428 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 25750 179200 25862 180000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 153262 179200 153374 180000 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 0 123708 800 123948 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 165498 179200 165610 180000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 86286 179200 86398 180000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 136518 0 136630 800 6 io_in[27]
port 21 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 117198 0 117310 800 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 35410 179200 35522 180000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 7074 179200 7186 180000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 48290 179200 48402 180000 6 io_in[31]
port 26 nsew signal input
rlabel metal3 s 0 73388 800 73628 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 179200 6748 180000 6988 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 94658 0 94770 800 6 io_in[34]
port 29 nsew signal input
rlabel metal3 s 179200 60468 180000 60708 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 0 163828 800 164068 6 io_in[36]
port 31 nsew signal input
rlabel metal3 s 179200 120988 180000 121228 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 151974 0 152086 800 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 0 147508 800 147748 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 59882 0 59994 800 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 79202 0 79314 800 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 148754 0 148866 800 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 0 16268 800 16508 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 120418 0 120530 800 6 io_oeb[0]
port 40 nsew signal bidirectional
rlabel metal2 s 130722 179200 130834 180000 6 io_oeb[10]
port 41 nsew signal bidirectional
rlabel metal2 s 158414 0 158526 800 6 io_oeb[11]
port 42 nsew signal bidirectional
rlabel metal2 s 137162 179200 137274 180000 6 io_oeb[12]
port 43 nsew signal bidirectional
rlabel metal3 s 179200 107388 180000 107628 6 io_oeb[13]
port 44 nsew signal bidirectional
rlabel metal3 s 179200 144788 180000 145028 6 io_oeb[14]
port 45 nsew signal bidirectional
rlabel metal3 s 179200 104668 180000 104908 6 io_oeb[15]
port 46 nsew signal bidirectional
rlabel metal3 s 0 59788 800 60028 6 io_oeb[16]
port 47 nsew signal bidirectional
rlabel metal2 s 88862 0 88974 800 6 io_oeb[17]
port 48 nsew signal bidirectional
rlabel metal2 s 162278 179200 162390 180000 6 io_oeb[18]
port 49 nsew signal bidirectional
rlabel metal3 s 0 33268 800 33508 6 io_oeb[19]
port 50 nsew signal bidirectional
rlabel metal3 s 179200 10148 180000 10388 6 io_oeb[1]
port 51 nsew signal bidirectional
rlabel metal3 s 0 2668 800 2908 6 io_oeb[20]
port 52 nsew signal bidirectional
rlabel metal2 s 50222 0 50334 800 6 io_oeb[21]
port 53 nsew signal bidirectional
rlabel metal3 s 179200 164508 180000 164748 6 io_oeb[22]
port 54 nsew signal bidirectional
rlabel metal2 s 146822 179200 146934 180000 6 io_oeb[23]
port 55 nsew signal bidirectional
rlabel metal2 s 15446 0 15558 800 6 io_oeb[24]
port 56 nsew signal bidirectional
rlabel metal2 s 56662 0 56774 800 6 io_oeb[25]
port 57 nsew signal bidirectional
rlabel metal3 s 179200 101268 180000 101508 6 io_oeb[26]
port 58 nsew signal bidirectional
rlabel metal2 s 113978 0 114090 800 6 io_oeb[27]
port 59 nsew signal bidirectional
rlabel metal3 s 0 56388 800 56628 6 io_oeb[28]
port 60 nsew signal bidirectional
rlabel metal2 s 83066 179200 83178 180000 6 io_oeb[29]
port 61 nsew signal bidirectional
rlabel metal3 s 0 133908 800 134148 6 io_oeb[2]
port 62 nsew signal bidirectional
rlabel metal2 s 16090 179200 16202 180000 6 io_oeb[30]
port 63 nsew signal bidirectional
rlabel metal2 s 175158 179200 175270 180000 6 io_oeb[31]
port 64 nsew signal bidirectional
rlabel metal2 s 102386 179200 102498 180000 6 io_oeb[32]
port 65 nsew signal bidirectional
rlabel metal3 s 179200 154988 180000 155228 6 io_oeb[33]
port 66 nsew signal bidirectional
rlabel metal3 s 179200 157708 180000 157948 6 io_oeb[34]
port 67 nsew signal bidirectional
rlabel metal3 s 0 90388 800 90628 6 io_oeb[35]
port 68 nsew signal bidirectional
rlabel metal2 s 150042 179200 150154 180000 6 io_oeb[36]
port 69 nsew signal bidirectional
rlabel metal3 s 179200 114188 180000 114428 6 io_oeb[37]
port 70 nsew signal bidirectional
rlabel metal2 s 32190 179200 32302 180000 6 io_oeb[3]
port 71 nsew signal bidirectional
rlabel metal3 s 179200 50948 180000 51188 6 io_oeb[4]
port 72 nsew signal bidirectional
rlabel metal3 s 0 150228 800 150468 6 io_oeb[5]
port 73 nsew signal bidirectional
rlabel metal2 s 19310 179200 19422 180000 6 io_oeb[6]
port 74 nsew signal bidirectional
rlabel metal3 s 179200 167908 180000 168148 6 io_oeb[7]
port 75 nsew signal bidirectional
rlabel metal3 s 179200 87668 180000 87908 6 io_oeb[8]
port 76 nsew signal bidirectional
rlabel metal3 s 0 76788 800 77028 6 io_oeb[9]
port 77 nsew signal bidirectional
rlabel metal3 s 0 170628 800 170868 6 io_out[0]
port 78 nsew signal bidirectional
rlabel metal3 s 0 6068 800 6308 6 io_out[10]
port 79 nsew signal bidirectional
rlabel metal2 s 97878 0 97990 800 6 io_out[11]
port 80 nsew signal bidirectional
rlabel metal3 s 0 80188 800 80428 6 io_out[12]
port 81 nsew signal bidirectional
rlabel metal2 s 111402 179200 111514 180000 6 io_out[13]
port 82 nsew signal bidirectional
rlabel metal2 s 178378 179200 178490 180000 6 io_out[14]
port 83 nsew signal bidirectional
rlabel metal3 s 0 120308 800 120548 6 io_out[15]
port 84 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 io_out[16]
port 85 nsew signal bidirectional
rlabel metal2 s 66966 179200 67078 180000 6 io_out[17]
port 86 nsew signal bidirectional
rlabel metal3 s 179200 40748 180000 40988 6 io_out[18]
port 87 nsew signal bidirectional
rlabel metal2 s 156482 179200 156594 180000 6 io_out[19]
port 88 nsew signal bidirectional
rlabel metal3 s 0 9468 800 9708 6 io_out[1]
port 89 nsew signal bidirectional
rlabel metal3 s 0 66588 800 66828 6 io_out[20]
port 90 nsew signal bidirectional
rlabel metal2 s 155194 0 155306 800 6 io_out[21]
port 91 nsew signal bidirectional
rlabel metal2 s 171938 179200 172050 180000 6 io_out[22]
port 92 nsew signal bidirectional
rlabel metal2 s 121062 179200 121174 180000 6 io_out[23]
port 93 nsew signal bidirectional
rlabel metal3 s 179200 110788 180000 111028 6 io_out[24]
port 94 nsew signal bidirectional
rlabel metal3 s 0 137308 800 137548 6 io_out[25]
port 95 nsew signal bidirectional
rlabel metal2 s 177734 0 177846 800 6 io_out[26]
port 96 nsew signal bidirectional
rlabel metal3 s 179200 77468 180000 77708 6 io_out[27]
port 97 nsew signal bidirectional
rlabel metal2 s 108826 179200 108938 180000 6 io_out[28]
port 98 nsew signal bidirectional
rlabel metal2 s 133942 179200 134054 180000 6 io_out[29]
port 99 nsew signal bidirectional
rlabel metal3 s 179200 57068 180000 57308 6 io_out[2]
port 100 nsew signal bidirectional
rlabel metal3 s 0 12868 800 13108 6 io_out[30]
port 101 nsew signal bidirectional
rlabel metal2 s 117842 179200 117954 180000 6 io_out[31]
port 102 nsew signal bidirectional
rlabel metal2 s 45070 179200 45182 180000 6 io_out[32]
port 103 nsew signal bidirectional
rlabel metal2 s 73406 179200 73518 180000 6 io_out[33]
port 104 nsew signal bidirectional
rlabel metal2 s 99166 179200 99278 180000 6 io_out[34]
port 105 nsew signal bidirectional
rlabel metal2 s 174514 0 174626 800 6 io_out[35]
port 106 nsew signal bidirectional
rlabel metal3 s 0 40068 800 40308 6 io_out[36]
port 107 nsew signal bidirectional
rlabel metal3 s 179200 13548 180000 13788 6 io_out[37]
port 108 nsew signal bidirectional
rlabel metal2 s 28326 0 28438 800 6 io_out[3]
port 109 nsew signal bidirectional
rlabel metal3 s 0 99908 800 100148 6 io_out[4]
port 110 nsew signal bidirectional
rlabel metal2 s 95946 179200 96058 180000 6 io_out[5]
port 111 nsew signal bidirectional
rlabel metal3 s 179200 80868 180000 81108 6 io_out[6]
port 112 nsew signal bidirectional
rlabel metal3 s 179200 33948 180000 34188 6 io_out[7]
port 113 nsew signal bidirectional
rlabel metal3 s 0 174028 800 174268 6 io_out[8]
port 114 nsew signal bidirectional
rlabel metal3 s 179200 151588 180000 151828 6 io_out[9]
port 115 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 117 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 117 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 117 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 117 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 117 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 117 nsew ground bidirectional
rlabel metal2 s 61170 179200 61282 180000 6 wb_clk_i
port 118 nsew signal input
rlabel metal3 s 179200 174708 180000 174948 6 wb_rst_i
port 119 nsew signal input
rlabel metal3 s 0 130508 800 130748 6 wbs_ack_o
port 120 nsew signal bidirectional
rlabel metal3 s 179200 117588 180000 117828 6 wbs_adr_i[0]
port 121 nsew signal input
rlabel metal3 s 179200 148188 180000 148428 6 wbs_adr_i[10]
port 122 nsew signal input
rlabel metal3 s 0 106708 800 106948 6 wbs_adr_i[11]
port 123 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 wbs_adr_i[12]
port 124 nsew signal input
rlabel metal2 s 69542 0 69654 800 6 wbs_adr_i[13]
port 125 nsew signal input
rlabel metal3 s 179200 44148 180000 44388 6 wbs_adr_i[14]
port 126 nsew signal input
rlabel metal2 s 92726 179200 92838 180000 6 wbs_adr_i[15]
port 127 nsew signal input
rlabel metal2 s 82422 0 82534 800 6 wbs_adr_i[16]
port 128 nsew signal input
rlabel metal3 s 179200 30548 180000 30788 6 wbs_adr_i[17]
port 129 nsew signal input
rlabel metal2 s 171294 0 171406 800 6 wbs_adr_i[18]
port 130 nsew signal input
rlabel metal3 s 0 160428 800 160668 6 wbs_adr_i[19]
port 131 nsew signal input
rlabel metal3 s 0 116908 800 117148 6 wbs_adr_i[1]
port 132 nsew signal input
rlabel metal3 s 179200 97868 180000 98108 6 wbs_adr_i[20]
port 133 nsew signal input
rlabel metal3 s 0 144108 800 144348 6 wbs_adr_i[21]
port 134 nsew signal input
rlabel metal3 s 0 63188 800 63428 6 wbs_adr_i[22]
port 135 nsew signal input
rlabel metal2 s 164854 0 164966 800 6 wbs_adr_i[23]
port 136 nsew signal input
rlabel metal2 s 54730 179200 54842 180000 6 wbs_adr_i[24]
port 137 nsew signal input
rlabel metal2 s 72762 0 72874 800 6 wbs_adr_i[25]
port 138 nsew signal input
rlabel metal3 s 0 86988 800 87228 6 wbs_adr_i[26]
port 139 nsew signal input
rlabel metal3 s 0 113508 800 113748 6 wbs_adr_i[27]
port 140 nsew signal input
rlabel metal3 s 0 52988 800 53228 6 wbs_adr_i[28]
port 141 nsew signal input
rlabel metal2 s 51510 179200 51622 180000 6 wbs_adr_i[29]
port 142 nsew signal input
rlabel metal2 s 53442 0 53554 800 6 wbs_adr_i[2]
port 143 nsew signal input
rlabel metal2 s 22530 179200 22642 180000 6 wbs_adr_i[30]
port 144 nsew signal input
rlabel metal3 s 179200 16948 180000 17188 6 wbs_adr_i[31]
port 145 nsew signal input
rlabel metal2 s 107538 0 107650 800 6 wbs_adr_i[3]
port 146 nsew signal input
rlabel metal3 s 179200 141388 180000 141628 6 wbs_adr_i[4]
port 147 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 wbs_adr_i[5]
port 148 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 wbs_adr_i[6]
port 149 nsew signal input
rlabel metal2 s 38630 179200 38742 180000 6 wbs_adr_i[7]
port 150 nsew signal input
rlabel metal2 s 142314 0 142426 800 6 wbs_adr_i[8]
port 151 nsew signal input
rlabel metal3 s 0 110108 800 110348 6 wbs_adr_i[9]
port 152 nsew signal input
rlabel metal2 s 143602 179200 143714 180000 6 wbs_cyc_i
port 153 nsew signal input
rlabel metal2 s 3854 179200 3966 180000 6 wbs_dat_i[0]
port 154 nsew signal input
rlabel metal2 s 41850 179200 41962 180000 6 wbs_dat_i[10]
port 155 nsew signal input
rlabel metal2 s 70186 179200 70298 180000 6 wbs_dat_i[11]
port 156 nsew signal input
rlabel metal2 s 63746 179200 63858 180000 6 wbs_dat_i[12]
port 157 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 wbs_dat_i[13]
port 158 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 wbs_dat_i[14]
port 159 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 wbs_dat_i[15]
port 160 nsew signal input
rlabel metal2 s 85642 0 85754 800 6 wbs_dat_i[16]
port 161 nsew signal input
rlabel metal3 s 179200 171308 180000 171548 6 wbs_dat_i[17]
port 162 nsew signal input
rlabel metal2 s 10294 179200 10406 180000 6 wbs_dat_i[18]
port 163 nsew signal input
rlabel metal2 s 89506 179200 89618 180000 6 wbs_dat_i[19]
port 164 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 wbs_dat_i[1]
port 165 nsew signal input
rlabel metal3 s 179200 63868 180000 64108 6 wbs_dat_i[20]
port 166 nsew signal input
rlabel metal3 s 179200 134588 180000 134828 6 wbs_dat_i[21]
port 167 nsew signal input
rlabel metal3 s 0 83588 800 83828 6 wbs_dat_i[22]
port 168 nsew signal input
rlabel metal3 s 179200 94468 180000 94708 6 wbs_dat_i[23]
port 169 nsew signal input
rlabel metal3 s 0 157028 800 157268 6 wbs_dat_i[24]
port 170 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 wbs_dat_i[25]
port 171 nsew signal input
rlabel metal3 s 179200 161108 180000 161348 6 wbs_dat_i[26]
port 172 nsew signal input
rlabel metal2 s 105606 179200 105718 180000 6 wbs_dat_i[27]
port 173 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 wbs_dat_i[28]
port 174 nsew signal input
rlabel metal3 s 179200 70668 180000 70908 6 wbs_dat_i[29]
port 175 nsew signal input
rlabel metal2 s 126858 0 126970 800 6 wbs_dat_i[2]
port 176 nsew signal input
rlabel metal3 s 179200 23748 180000 23988 6 wbs_dat_i[30]
port 177 nsew signal input
rlabel metal3 s 0 167228 800 167468 6 wbs_dat_i[31]
port 178 nsew signal input
rlabel metal2 s 161634 0 161746 800 6 wbs_dat_i[3]
port 179 nsew signal input
rlabel metal2 s 25106 0 25218 800 6 wbs_dat_i[4]
port 180 nsew signal input
rlabel metal2 s 75982 0 76094 800 6 wbs_dat_i[5]
port 181 nsew signal input
rlabel metal3 s 179200 47548 180000 47788 6 wbs_dat_i[6]
port 182 nsew signal input
rlabel metal3 s 179200 178108 180000 178348 6 wbs_dat_i[7]
port 183 nsew signal input
rlabel metal3 s 0 46868 800 47108 6 wbs_dat_i[8]
port 184 nsew signal input
rlabel metal2 s 168074 0 168186 800 6 wbs_dat_i[9]
port 185 nsew signal input
rlabel metal3 s 0 69988 800 70228 6 wbs_dat_o[0]
port 186 nsew signal bidirectional
rlabel metal3 s 179200 74068 180000 74308 6 wbs_dat_o[10]
port 187 nsew signal bidirectional
rlabel metal2 s 2566 0 2678 800 6 wbs_dat_o[11]
port 188 nsew signal bidirectional
rlabel metal3 s 179200 137988 180000 138228 6 wbs_dat_o[12]
port 189 nsew signal bidirectional
rlabel metal2 s 168718 179200 168830 180000 6 wbs_dat_o[13]
port 190 nsew signal bidirectional
rlabel metal3 s 179200 628 180000 868 6 wbs_dat_o[14]
port 191 nsew signal bidirectional
rlabel metal2 s 159058 179200 159170 180000 6 wbs_dat_o[15]
port 192 nsew signal bidirectional
rlabel metal3 s 0 97188 800 97428 6 wbs_dat_o[16]
port 193 nsew signal bidirectional
rlabel metal3 s 0 103308 800 103548 6 wbs_dat_o[17]
port 194 nsew signal bidirectional
rlabel metal2 s 110758 0 110870 800 6 wbs_dat_o[18]
port 195 nsew signal bidirectional
rlabel metal2 s -10 0 102 800 6 wbs_dat_o[19]
port 196 nsew signal bidirectional
rlabel metal2 s 130078 0 130190 800 6 wbs_dat_o[1]
port 197 nsew signal bidirectional
rlabel metal3 s 0 127108 800 127348 6 wbs_dat_o[20]
port 198 nsew signal bidirectional
rlabel metal2 s 13514 179200 13626 180000 6 wbs_dat_o[21]
port 199 nsew signal bidirectional
rlabel metal2 s 79846 179200 79958 180000 6 wbs_dat_o[22]
port 200 nsew signal bidirectional
rlabel metal3 s 0 93788 800 94028 6 wbs_dat_o[23]
port 201 nsew signal bidirectional
rlabel metal2 s 34766 0 34878 800 6 wbs_dat_o[24]
port 202 nsew signal bidirectional
rlabel metal2 s 12226 0 12338 800 6 wbs_dat_o[25]
port 203 nsew signal bidirectional
rlabel metal2 s 114622 179200 114734 180000 6 wbs_dat_o[26]
port 204 nsew signal bidirectional
rlabel metal2 s 76626 179200 76738 180000 6 wbs_dat_o[27]
port 205 nsew signal bidirectional
rlabel metal2 s 92082 0 92194 800 6 wbs_dat_o[28]
port 206 nsew signal bidirectional
rlabel metal2 s 140382 179200 140494 180000 6 wbs_dat_o[29]
port 207 nsew signal bidirectional
rlabel metal3 s 179200 37348 180000 37588 6 wbs_dat_o[2]
port 208 nsew signal bidirectional
rlabel metal3 s 0 140708 800 140948 6 wbs_dat_o[30]
port 209 nsew signal bidirectional
rlabel metal3 s 179200 127788 180000 128028 6 wbs_dat_o[31]
port 210 nsew signal bidirectional
rlabel metal2 s 37986 0 38098 800 6 wbs_dat_o[3]
port 211 nsew signal bidirectional
rlabel metal2 s 63102 0 63214 800 6 wbs_dat_o[4]
port 212 nsew signal bidirectional
rlabel metal2 s 101098 0 101210 800 6 wbs_dat_o[5]
port 213 nsew signal bidirectional
rlabel metal3 s 179200 124388 180000 124628 6 wbs_dat_o[6]
port 214 nsew signal bidirectional
rlabel metal2 s 104318 0 104430 800 6 wbs_dat_o[7]
port 215 nsew signal bidirectional
rlabel metal2 s 127502 179200 127614 180000 6 wbs_dat_o[8]
port 216 nsew signal bidirectional
rlabel metal2 s 124282 179200 124394 180000 6 wbs_dat_o[9]
port 217 nsew signal bidirectional
rlabel metal3 s 0 177428 800 177668 6 wbs_sel_i[0]
port 218 nsew signal input
rlabel metal2 s 28970 179200 29082 180000 6 wbs_sel_i[1]
port 219 nsew signal input
rlabel metal2 s 123638 0 123750 800 6 wbs_sel_i[2]
port 220 nsew signal input
rlabel metal3 s 0 43468 800 43708 6 wbs_sel_i[3]
port 221 nsew signal input
rlabel metal3 s 0 153628 800 153868 6 wbs_stb_i
port 222 nsew signal input
rlabel metal3 s 179200 84268 180000 84508 6 wbs_we_i
port 223 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 32254634
string GDS_FILE /home/runner/caravel_user_project/openlane/wrapped_etpu/runs/22_08_28_18_54/results/signoff/wrapped_etpu.magic.gds
string GDS_START 891348
<< end >>

