magic
tech sky130B
magscale 1 2
timestamp 1660477629
<< viali >>
rect 67465 69445 67499 69479
rect 1501 69377 1535 69411
rect 55505 69377 55539 69411
rect 2053 69309 2087 69343
rect 55781 69309 55815 69343
rect 67649 69241 67683 69275
rect 46765 69173 46799 69207
rect 51273 69173 51307 69207
rect 56977 69173 57011 69207
rect 59277 69173 59311 69207
rect 46489 68833 46523 68867
rect 46949 68833 46983 68867
rect 50997 68833 51031 68867
rect 51549 68833 51583 68867
rect 56241 68833 56275 68867
rect 57069 68833 57103 68867
rect 48789 68765 48823 68799
rect 58909 68765 58943 68799
rect 46673 68697 46707 68731
rect 51181 68697 51215 68731
rect 56425 68697 56459 68731
rect 48881 68629 48915 68663
rect 59001 68629 59035 68663
rect 51181 68425 51215 68459
rect 56425 68425 56459 68459
rect 51089 68289 51123 68323
rect 56333 68289 56367 68323
rect 59001 68289 59035 68323
rect 59185 68221 59219 68255
rect 60841 68221 60875 68255
rect 60933 67677 60967 67711
rect 61117 67609 61151 67643
rect 62773 67609 62807 67643
rect 60657 67337 60691 67371
rect 60565 67201 60599 67235
rect 61393 67201 61427 67235
rect 37749 66589 37783 66623
rect 44097 66589 44131 66623
rect 37473 66113 37507 66147
rect 43821 66113 43855 66147
rect 37657 66045 37691 66079
rect 38669 66045 38703 66079
rect 44005 66045 44039 66079
rect 45477 66045 45511 66079
rect 37749 65705 37783 65739
rect 43821 65705 43855 65739
rect 7021 65501 7055 65535
rect 31861 65501 31895 65535
rect 32321 65501 32355 65535
rect 37657 65501 37691 65535
rect 42901 65501 42935 65535
rect 43729 65501 43763 65535
rect 32597 65433 32631 65467
rect 31493 65093 31527 65127
rect 32321 65093 32355 65127
rect 6745 65025 6779 65059
rect 31401 65025 31435 65059
rect 42625 65025 42659 65059
rect 6929 64957 6963 64991
rect 7205 64957 7239 64991
rect 30941 64957 30975 64991
rect 32137 64957 32171 64991
rect 33149 64957 33183 64991
rect 42809 64957 42843 64991
rect 44189 64957 44223 64991
rect 55965 64821 55999 64855
rect 7113 64617 7147 64651
rect 30481 64617 30515 64651
rect 30941 64617 30975 64651
rect 42809 64617 42843 64651
rect 31033 64549 31067 64583
rect 31217 64549 31251 64583
rect 31677 64481 31711 64515
rect 32137 64481 32171 64515
rect 55689 64481 55723 64515
rect 57529 64481 57563 64515
rect 7021 64413 7055 64447
rect 29745 64413 29779 64447
rect 30205 64413 30239 64447
rect 33977 64413 34011 64447
rect 34161 64413 34195 64447
rect 42717 64413 42751 64447
rect 30849 64345 30883 64379
rect 31217 64345 31251 64379
rect 31861 64345 31895 64379
rect 55873 64345 55907 64379
rect 34069 64277 34103 64311
rect 55689 64073 55723 64107
rect 28733 64005 28767 64039
rect 29469 64005 29503 64039
rect 31125 64005 31159 64039
rect 33977 64005 34011 64039
rect 28641 63937 28675 63971
rect 32137 63937 32171 63971
rect 55597 63937 55631 63971
rect 29285 63869 29319 63903
rect 32321 63869 32355 63903
rect 58081 63733 58115 63767
rect 33241 63461 33275 63495
rect 31309 63393 31343 63427
rect 57621 63393 57655 63427
rect 59093 63393 59127 63427
rect 30665 63325 30699 63359
rect 31565 63325 31599 63359
rect 33149 63325 33183 63359
rect 50353 63325 50387 63359
rect 30757 63257 30791 63291
rect 57805 63257 57839 63291
rect 32689 63189 32723 63223
rect 49157 62985 49191 63019
rect 57989 62985 58023 63019
rect 48973 62849 49007 62883
rect 49709 62849 49743 62883
rect 57897 62849 57931 62883
rect 64981 62849 65015 62883
rect 31585 62781 31619 62815
rect 32137 62781 32171 62815
rect 32321 62781 32355 62815
rect 32597 62781 32631 62815
rect 49893 62781 49927 62815
rect 50353 62781 50387 62815
rect 65809 62713 65843 62747
rect 46765 62645 46799 62679
rect 65073 62645 65107 62679
rect 32413 62441 32447 62475
rect 50261 62441 50295 62475
rect 46489 62305 46523 62339
rect 48237 62305 48271 62339
rect 67465 62305 67499 62339
rect 32321 62237 32355 62271
rect 50169 62237 50203 62271
rect 54677 62237 54711 62271
rect 65073 62237 65107 62271
rect 65625 62237 65659 62271
rect 46673 62169 46707 62203
rect 65809 62169 65843 62203
rect 46673 61897 46707 61931
rect 64613 61897 64647 61931
rect 65349 61829 65383 61863
rect 67005 61829 67039 61863
rect 46581 61761 46615 61795
rect 54493 61761 54527 61795
rect 64521 61761 64555 61795
rect 65165 61761 65199 61795
rect 54677 61693 54711 61727
rect 56333 61693 56367 61727
rect 54493 61353 54527 61387
rect 23213 61149 23247 61183
rect 54401 61149 54435 61183
rect 23029 60673 23063 60707
rect 1409 60605 1443 60639
rect 1685 60605 1719 60639
rect 23213 60605 23247 60639
rect 23673 60605 23707 60639
rect 23581 60265 23615 60299
rect 47593 60129 47627 60163
rect 23489 60061 23523 60095
rect 26985 60061 27019 60095
rect 46673 60061 46707 60095
rect 47133 60061 47167 60095
rect 47317 59993 47351 60027
rect 47685 59721 47719 59755
rect 28825 59653 28859 59687
rect 47593 59585 47627 59619
rect 26433 59517 26467 59551
rect 26985 59517 27019 59551
rect 27169 59517 27203 59551
rect 26249 59177 26283 59211
rect 26801 59041 26835 59075
rect 27261 59041 27295 59075
rect 26157 58973 26191 59007
rect 26985 58905 27019 58939
rect 27169 58633 27203 58667
rect 27077 58497 27111 58531
rect 48697 57885 48731 57919
rect 48421 57409 48455 57443
rect 48605 57341 48639 57375
rect 48881 57341 48915 57375
rect 48605 57001 48639 57035
rect 11621 56865 11655 56899
rect 10701 56797 10735 56831
rect 11161 56797 11195 56831
rect 48513 56797 48547 56831
rect 11345 56729 11379 56763
rect 11621 56457 11655 56491
rect 11529 56321 11563 56355
rect 57345 55709 57379 55743
rect 32781 55301 32815 55335
rect 37381 55301 37415 55335
rect 57069 55301 57103 55335
rect 58081 55301 58115 55335
rect 32597 55233 32631 55267
rect 37289 55233 37323 55267
rect 56977 55233 57011 55267
rect 57897 55233 57931 55267
rect 59737 55233 59771 55267
rect 33057 55165 33091 55199
rect 27537 53941 27571 53975
rect 39037 53941 39071 53975
rect 51457 53941 51491 53975
rect 67649 53941 67683 53975
rect 27169 53601 27203 53635
rect 27629 53601 27663 53635
rect 51181 53601 51215 53635
rect 66269 53601 66303 53635
rect 66729 53601 66763 53635
rect 27353 53465 27387 53499
rect 51365 53465 51399 53499
rect 53021 53465 53055 53499
rect 66453 53465 66487 53499
rect 27905 53193 27939 53227
rect 51181 53193 51215 53227
rect 67557 53193 67591 53227
rect 38301 53125 38335 53159
rect 39037 53125 39071 53159
rect 40693 53125 40727 53159
rect 27813 53057 27847 53091
rect 38209 53057 38243 53091
rect 38853 53057 38887 53091
rect 51089 53057 51123 53091
rect 67465 53057 67499 53091
rect 5549 52853 5583 52887
rect 7849 52853 7883 52887
rect 5273 52513 5307 52547
rect 5457 52513 5491 52547
rect 5733 52513 5767 52547
rect 8125 52445 8159 52479
rect 8217 52309 8251 52343
rect 5733 52105 5767 52139
rect 7757 52037 7791 52071
rect 5641 51969 5675 52003
rect 7573 51969 7607 52003
rect 8033 51901 8067 51935
rect 51641 51765 51675 51799
rect 51365 51425 51399 51459
rect 53205 51425 53239 51459
rect 35541 51357 35575 51391
rect 45569 51357 45603 51391
rect 51549 51289 51583 51323
rect 51365 51017 51399 51051
rect 36737 50949 36771 50983
rect 34897 50881 34931 50915
rect 45201 50881 45235 50915
rect 51273 50881 51307 50915
rect 35081 50813 35115 50847
rect 45385 50813 45419 50847
rect 45661 50813 45695 50847
rect 63693 50677 63727 50711
rect 35357 50473 35391 50507
rect 46029 50473 46063 50507
rect 63233 50337 63267 50371
rect 64797 50337 64831 50371
rect 7205 50269 7239 50303
rect 28733 50269 28767 50303
rect 30297 50269 30331 50303
rect 35265 50269 35299 50303
rect 45937 50269 45971 50303
rect 63417 50201 63451 50235
rect 63233 49929 63267 49963
rect 29285 49861 29319 49895
rect 6929 49793 6963 49827
rect 27445 49793 27479 49827
rect 29745 49793 29779 49827
rect 63141 49793 63175 49827
rect 7113 49725 7147 49759
rect 7389 49725 7423 49759
rect 27629 49725 27663 49759
rect 29929 49725 29963 49759
rect 31125 49725 31159 49759
rect 7297 49385 7331 49419
rect 28641 49385 28675 49419
rect 30389 49385 30423 49419
rect 7205 49181 7239 49215
rect 28549 49181 28583 49215
rect 30297 49181 30331 49215
rect 54125 49181 54159 49215
rect 44465 48773 44499 48807
rect 53297 48773 53331 48807
rect 54033 48773 54067 48807
rect 55689 48773 55723 48807
rect 43545 48705 43579 48739
rect 44189 48705 44223 48739
rect 45201 48705 45235 48739
rect 53205 48705 53239 48739
rect 53849 48705 53883 48739
rect 45477 48637 45511 48671
rect 43637 48501 43671 48535
rect 44005 48229 44039 48263
rect 43269 48093 43303 48127
rect 45017 48093 45051 48127
rect 43821 48025 43855 48059
rect 45293 48025 45327 48059
rect 43637 47685 43671 47719
rect 64797 47685 64831 47719
rect 65533 47685 65567 47719
rect 43453 47617 43487 47651
rect 64705 47617 64739 47651
rect 43913 47549 43947 47583
rect 65349 47549 65383 47583
rect 67189 47549 67223 47583
rect 65809 47209 65843 47243
rect 43637 47073 43671 47107
rect 43913 47073 43947 47107
rect 45385 47073 45419 47107
rect 45109 47005 45143 47039
rect 37381 45917 37415 45951
rect 37289 45441 37323 45475
rect 49525 45441 49559 45475
rect 37473 45373 37507 45407
rect 38485 45373 38519 45407
rect 49801 45305 49835 45339
rect 14933 45237 14967 45271
rect 67649 45237 67683 45271
rect 36921 45033 36955 45067
rect 14749 44897 14783 44931
rect 15209 44897 15243 44931
rect 66269 44897 66303 44931
rect 68109 44897 68143 44931
rect 36829 44829 36863 44863
rect 14933 44761 14967 44795
rect 66453 44761 66487 44795
rect 15117 44489 15151 44523
rect 67557 44489 67591 44523
rect 15025 44353 15059 44387
rect 37749 44353 37783 44387
rect 44097 44353 44131 44387
rect 67465 44353 67499 44387
rect 38025 44285 38059 44319
rect 44189 44149 44223 44183
rect 52101 43741 52135 43775
rect 52745 43741 52779 43775
rect 52193 43673 52227 43707
rect 52929 43673 52963 43707
rect 54585 43673 54619 43707
rect 53021 43265 53055 43299
rect 54493 42653 54527 42687
rect 54585 42517 54619 42551
rect 54953 42245 54987 42279
rect 19993 42177 20027 42211
rect 44097 42177 44131 42211
rect 20821 42109 20855 42143
rect 44281 42109 44315 42143
rect 54309 42109 54343 42143
rect 54769 42109 54803 42143
rect 56517 42109 56551 42143
rect 57253 41157 57287 41191
rect 58081 41157 58115 41191
rect 57161 41089 57195 41123
rect 57897 41021 57931 41055
rect 59737 41021 59771 41055
rect 57897 40681 57931 40715
rect 9781 39797 9815 39831
rect 35357 39797 35391 39831
rect 60749 39797 60783 39831
rect 63877 39797 63911 39831
rect 9597 39457 9631 39491
rect 10057 39457 10091 39491
rect 23121 39457 23155 39491
rect 35081 39457 35115 39491
rect 36921 39457 36955 39491
rect 60473 39457 60507 39491
rect 62037 39457 62071 39491
rect 63233 39457 63267 39491
rect 64797 39457 64831 39491
rect 22477 39389 22511 39423
rect 9781 39321 9815 39355
rect 35265 39321 35299 39355
rect 60657 39321 60691 39355
rect 63417 39321 63451 39355
rect 9873 39049 9907 39083
rect 34897 39049 34931 39083
rect 60473 39049 60507 39083
rect 63509 39049 63543 39083
rect 24133 38981 24167 39015
rect 9781 38913 9815 38947
rect 22293 38913 22327 38947
rect 34805 38913 34839 38947
rect 44649 38913 44683 38947
rect 47685 38913 47719 38947
rect 47961 38913 47995 38947
rect 60381 38913 60415 38947
rect 63417 38913 63451 38947
rect 22477 38845 22511 38879
rect 44741 38709 44775 38743
rect 21465 38505 21499 38539
rect 32781 38369 32815 38403
rect 45201 38369 45235 38403
rect 21373 38301 21407 38335
rect 22017 38301 22051 38335
rect 23857 38301 23891 38335
rect 32321 38301 32355 38335
rect 44465 38301 44499 38335
rect 45017 38301 45051 38335
rect 51549 38301 51583 38335
rect 22201 38233 22235 38267
rect 32505 38233 32539 38267
rect 46857 38233 46891 38267
rect 22661 37961 22695 37995
rect 33517 37961 33551 37995
rect 20821 37893 20855 37927
rect 6653 37825 6687 37859
rect 20545 37825 20579 37859
rect 22569 37825 22603 37859
rect 32965 37825 32999 37859
rect 33425 37825 33459 37859
rect 48789 37825 48823 37859
rect 51181 37825 51215 37859
rect 49065 37757 49099 37791
rect 6745 37621 6779 37655
rect 51273 37621 51307 37655
rect 20085 37281 20119 37315
rect 51365 37281 51399 37315
rect 5457 37213 5491 37247
rect 6469 37213 6503 37247
rect 19809 37213 19843 37247
rect 20637 37213 20671 37247
rect 21557 37213 21591 37247
rect 21833 37213 21867 37247
rect 53205 37213 53239 37247
rect 20913 37145 20947 37179
rect 51549 37145 51583 37179
rect 6561 36805 6595 36839
rect 5457 36737 5491 36771
rect 6377 36737 6411 36771
rect 20637 36737 20671 36771
rect 38853 36737 38887 36771
rect 6837 36669 6871 36703
rect 20913 36669 20947 36703
rect 5549 36533 5583 36567
rect 38393 36533 38427 36567
rect 38945 36533 38979 36567
rect 20545 36329 20579 36363
rect 5273 36193 5307 36227
rect 5457 36193 5491 36227
rect 5733 36193 5767 36227
rect 20729 36125 20763 36159
rect 38301 35717 38335 35751
rect 37381 35649 37415 35683
rect 38117 35649 38151 35683
rect 39773 35581 39807 35615
rect 63049 35581 63083 35615
rect 63233 35581 63267 35615
rect 64889 35581 64923 35615
rect 37473 35445 37507 35479
rect 63233 35241 63267 35275
rect 63785 35241 63819 35275
rect 37105 35105 37139 35139
rect 37381 35105 37415 35139
rect 36461 35037 36495 35071
rect 36921 35037 36955 35071
rect 63693 35037 63727 35071
rect 42441 33949 42475 33983
rect 43545 33949 43579 33983
rect 42717 33881 42751 33915
rect 41429 33473 41463 33507
rect 42901 33473 42935 33507
rect 67465 33473 67499 33507
rect 41613 33405 41647 33439
rect 43085 33405 43119 33439
rect 44741 33405 44775 33439
rect 62405 33269 62439 33303
rect 67557 33269 67591 33303
rect 43545 33065 43579 33099
rect 42165 32929 42199 32963
rect 62221 32929 62255 32963
rect 67925 32929 67959 32963
rect 42441 32861 42475 32895
rect 43453 32861 43487 32895
rect 44097 32861 44131 32895
rect 67097 32861 67131 32895
rect 62405 32793 62439 32827
rect 64061 32793 64095 32827
rect 44189 32725 44223 32759
rect 67189 32725 67223 32759
rect 61945 32521 61979 32555
rect 42717 32453 42751 32487
rect 44097 32453 44131 32487
rect 65993 32453 66027 32487
rect 42441 32385 42475 32419
rect 43913 32385 43947 32419
rect 61853 32385 61887 32419
rect 65809 32385 65843 32419
rect 45477 32317 45511 32351
rect 67557 32317 67591 32351
rect 66269 31841 66303 31875
rect 67833 31841 67867 31875
rect 42349 31773 42383 31807
rect 66453 31705 66487 31739
rect 42441 31637 42475 31671
rect 42625 31365 42659 31399
rect 59093 31365 59127 31399
rect 59829 31365 59863 31399
rect 59001 31297 59035 31331
rect 67649 31297 67683 31331
rect 41889 31229 41923 31263
rect 42441 31229 42475 31263
rect 42901 31229 42935 31263
rect 59645 31229 59679 31263
rect 61485 31229 61519 31263
rect 59829 30889 59863 30923
rect 26433 30685 26467 30719
rect 27077 30685 27111 30719
rect 42349 30685 42383 30719
rect 26525 30617 26559 30651
rect 27261 30617 27295 30651
rect 28917 30617 28951 30651
rect 42625 30617 42659 30651
rect 42901 30277 42935 30311
rect 27261 30209 27295 30243
rect 8033 30141 8067 30175
rect 8217 30141 8251 30175
rect 9137 30141 9171 30175
rect 42993 30005 43027 30039
rect 8217 29801 8251 29835
rect 9045 29801 9079 29835
rect 6101 29665 6135 29699
rect 4997 29597 5031 29631
rect 5641 29597 5675 29631
rect 8953 29597 8987 29631
rect 12449 29597 12483 29631
rect 43913 29597 43947 29631
rect 5089 29529 5123 29563
rect 5825 29529 5859 29563
rect 6561 29121 6595 29155
rect 12173 29121 12207 29155
rect 43637 29121 43671 29155
rect 12357 29053 12391 29087
rect 12817 29053 12851 29087
rect 43821 29053 43855 29087
rect 45201 29053 45235 29087
rect 12725 28713 12759 28747
rect 43637 28713 43671 28747
rect 4997 28509 5031 28543
rect 5457 28509 5491 28543
rect 12633 28509 12667 28543
rect 43545 28509 43579 28543
rect 54217 28509 54251 28543
rect 55321 28509 55355 28543
rect 54309 28441 54343 28475
rect 55505 28441 55539 28475
rect 57161 28441 57195 28475
rect 5549 28373 5583 28407
rect 9505 28033 9539 28067
rect 26985 28033 27019 28067
rect 54769 28033 54803 28067
rect 9597 27829 9631 27863
rect 10333 27829 10367 27863
rect 26249 27829 26283 27863
rect 27077 27829 27111 27863
rect 5089 27489 5123 27523
rect 5273 27489 5307 27523
rect 5641 27489 5675 27523
rect 9229 27489 9263 27523
rect 9413 27489 9447 27523
rect 9689 27489 9723 27523
rect 26065 27489 26099 27523
rect 26525 27489 26559 27523
rect 26249 27353 26283 27387
rect 34713 25857 34747 25891
rect 34805 25653 34839 25687
rect 35081 25313 35115 25347
rect 34897 25245 34931 25279
rect 36737 25177 36771 25211
rect 28825 24769 28859 24803
rect 35173 24769 35207 24803
rect 28365 24565 28399 24599
rect 28917 24565 28951 24599
rect 58449 24157 58483 24191
rect 28549 23749 28583 23783
rect 28365 23681 28399 23715
rect 58173 23681 58207 23715
rect 28825 23613 28859 23647
rect 58357 23613 58391 23647
rect 60013 23613 60047 23647
rect 57989 23273 58023 23307
rect 10793 23069 10827 23103
rect 11621 23069 11655 23103
rect 57897 23069 57931 23103
rect 60749 23069 60783 23103
rect 61577 23069 61611 23103
rect 10885 22933 10919 22967
rect 60841 22933 60875 22967
rect 60841 22661 60875 22695
rect 50537 22593 50571 22627
rect 60657 22593 60691 22627
rect 62497 22525 62531 22559
rect 4721 22389 4755 22423
rect 50629 22389 50663 22423
rect 51365 22389 51399 22423
rect 4537 22049 4571 22083
rect 4997 22049 5031 22083
rect 10793 22049 10827 22083
rect 12357 22049 12391 22083
rect 50537 22049 50571 22083
rect 50813 22049 50847 22083
rect 10609 21981 10643 22015
rect 50353 21981 50387 22015
rect 62957 21981 62991 22015
rect 4721 21913 4755 21947
rect 63049 21845 63083 21879
rect 5089 21641 5123 21675
rect 63325 21573 63359 21607
rect 4997 21505 5031 21539
rect 63141 21437 63175 21471
rect 64981 21437 65015 21471
rect 63325 21097 63359 21131
rect 32321 19805 32355 19839
rect 33977 19397 34011 19431
rect 32137 19329 32171 19363
rect 32321 19261 32355 19295
rect 32505 18921 32539 18955
rect 32413 18717 32447 18751
rect 5457 18037 5491 18071
rect 5181 17697 5215 17731
rect 6837 17697 6871 17731
rect 62681 17629 62715 17663
rect 63509 17629 63543 17663
rect 5365 17561 5399 17595
rect 62773 17493 62807 17527
rect 5549 17289 5583 17323
rect 63233 17221 63267 17255
rect 5457 17153 5491 17187
rect 63049 17153 63083 17187
rect 64797 17085 64831 17119
rect 13093 15453 13127 15487
rect 12817 14977 12851 15011
rect 13001 14909 13035 14943
rect 13553 14909 13587 14943
rect 12909 14569 12943 14603
rect 12817 14365 12851 14399
rect 19625 14365 19659 14399
rect 22109 14365 22143 14399
rect 22201 14229 22235 14263
rect 22201 13957 22235 13991
rect 19441 13889 19475 13923
rect 19625 13821 19659 13855
rect 19901 13821 19935 13855
rect 22017 13821 22051 13855
rect 22569 13821 22603 13855
rect 19993 13481 20027 13515
rect 22201 13481 22235 13515
rect 19901 13277 19935 13311
rect 35541 13277 35575 13311
rect 35633 13141 35667 13175
rect 35725 12597 35759 12631
rect 35449 12257 35483 12291
rect 35633 12257 35667 12291
rect 36093 12257 36127 12291
rect 34713 12189 34747 12223
rect 63601 12189 63635 12223
rect 34805 12053 34839 12087
rect 34437 11781 34471 11815
rect 63417 11713 63451 11747
rect 33793 11645 33827 11679
rect 34253 11645 34287 11679
rect 34805 11645 34839 11679
rect 63601 11645 63635 11679
rect 65257 11645 65291 11679
rect 24777 11509 24811 11543
rect 30297 11509 30331 11543
rect 63325 11305 63359 11339
rect 30573 11169 30607 11203
rect 35357 11169 35391 11203
rect 24593 11101 24627 11135
rect 26893 11101 26927 11135
rect 30113 11101 30147 11135
rect 34161 11101 34195 11135
rect 34897 11101 34931 11135
rect 63233 11101 63267 11135
rect 24777 11033 24811 11067
rect 26433 11033 26467 11067
rect 30297 11033 30331 11067
rect 35081 11033 35115 11067
rect 26985 10965 27019 10999
rect 25145 10761 25179 10795
rect 30665 10761 30699 10795
rect 35265 10761 35299 10795
rect 25053 10625 25087 10659
rect 30573 10625 30607 10659
rect 35173 10625 35207 10659
rect 26341 10421 26375 10455
rect 26065 10081 26099 10115
rect 26249 10081 26283 10115
rect 43361 10013 43395 10047
rect 27905 9945 27939 9979
rect 43453 9877 43487 9911
rect 43453 9605 43487 9639
rect 43269 9469 43303 9503
rect 43821 9469 43855 9503
rect 43545 9129 43579 9163
rect 26893 8993 26927 9027
rect 25973 8925 26007 8959
rect 26433 8925 26467 8959
rect 54401 8925 54435 8959
rect 55505 8925 55539 8959
rect 26617 8857 26651 8891
rect 54493 8789 54527 8823
rect 27077 8585 27111 8619
rect 54953 8517 54987 8551
rect 26985 8449 27019 8483
rect 54769 8449 54803 8483
rect 56609 8381 56643 8415
rect 27353 3553 27387 3587
rect 26893 3485 26927 3519
rect 40693 3485 40727 3519
rect 27077 3417 27111 3451
rect 40877 3417 40911 3451
rect 42533 3417 42567 3451
rect 41797 3145 41831 3179
rect 27077 3077 27111 3111
rect 27813 3077 27847 3111
rect 26433 3009 26467 3043
rect 26985 3009 27019 3043
rect 41705 3009 41739 3043
rect 27629 2941 27663 2975
rect 28089 2941 28123 2975
rect 38945 2941 38979 2975
rect 39405 2941 39439 2975
rect 39589 2941 39623 2975
rect 39957 2941 39991 2975
rect 27169 2601 27203 2635
rect 27905 2601 27939 2635
rect 39957 2601 39991 2635
rect 40877 2601 40911 2635
rect 27077 2397 27111 2431
rect 39865 2397 39899 2431
<< metal1 >>
rect 47394 71408 47400 71460
rect 47452 71448 47458 71460
rect 48222 71448 48228 71460
rect 47452 71420 48228 71448
rect 47452 71408 47458 71420
rect 48222 71408 48228 71420
rect 48280 71408 48286 71460
rect 1104 69658 68816 69680
rect 1104 69606 19574 69658
rect 19626 69606 19638 69658
rect 19690 69606 19702 69658
rect 19754 69606 19766 69658
rect 19818 69606 19830 69658
rect 19882 69606 50294 69658
rect 50346 69606 50358 69658
rect 50410 69606 50422 69658
rect 50474 69606 50486 69658
rect 50538 69606 50550 69658
rect 50602 69606 68816 69658
rect 1104 69584 68816 69606
rect 67450 69476 67456 69488
rect 67411 69448 67456 69476
rect 67450 69436 67456 69448
rect 67508 69436 67514 69488
rect 1486 69408 1492 69420
rect 1447 69380 1492 69408
rect 1486 69368 1492 69380
rect 1544 69368 1550 69420
rect 55398 69368 55404 69420
rect 55456 69408 55462 69420
rect 55493 69411 55551 69417
rect 55493 69408 55505 69411
rect 55456 69380 55505 69408
rect 55456 69368 55462 69380
rect 55493 69377 55505 69380
rect 55539 69377 55551 69411
rect 55493 69371 55551 69377
rect 2041 69343 2099 69349
rect 2041 69309 2053 69343
rect 2087 69340 2099 69343
rect 31386 69340 31392 69352
rect 2087 69312 31392 69340
rect 2087 69309 2099 69312
rect 2041 69303 2099 69309
rect 31386 69300 31392 69312
rect 31444 69300 31450 69352
rect 34054 69300 34060 69352
rect 34112 69340 34118 69352
rect 55769 69343 55827 69349
rect 55769 69340 55781 69343
rect 34112 69312 55781 69340
rect 34112 69300 34118 69312
rect 55769 69309 55781 69312
rect 55815 69309 55827 69343
rect 55769 69303 55827 69309
rect 30466 69232 30472 69284
rect 30524 69272 30530 69284
rect 67637 69275 67695 69281
rect 67637 69272 67649 69275
rect 30524 69244 67649 69272
rect 30524 69232 30530 69244
rect 67637 69241 67649 69244
rect 67683 69241 67695 69275
rect 67637 69235 67695 69241
rect 46750 69204 46756 69216
rect 46711 69176 46756 69204
rect 46750 69164 46756 69176
rect 46808 69164 46814 69216
rect 51258 69204 51264 69216
rect 51219 69176 51264 69204
rect 51258 69164 51264 69176
rect 51316 69164 51322 69216
rect 56962 69204 56968 69216
rect 56923 69176 56968 69204
rect 56962 69164 56968 69176
rect 57020 69164 57026 69216
rect 58986 69164 58992 69216
rect 59044 69204 59050 69216
rect 59265 69207 59323 69213
rect 59265 69204 59277 69207
rect 59044 69176 59277 69204
rect 59044 69164 59050 69176
rect 59265 69173 59277 69176
rect 59311 69173 59323 69207
rect 59265 69167 59323 69173
rect 1104 69114 68816 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 34934 69114
rect 34986 69062 34998 69114
rect 35050 69062 35062 69114
rect 35114 69062 35126 69114
rect 35178 69062 35190 69114
rect 35242 69062 65654 69114
rect 65706 69062 65718 69114
rect 65770 69062 65782 69114
rect 65834 69062 65846 69114
rect 65898 69062 65910 69114
rect 65962 69062 68816 69114
rect 1104 69040 68816 69062
rect 25130 68960 25136 69012
rect 25188 69000 25194 69012
rect 28258 69000 28264 69012
rect 25188 68972 28264 69000
rect 25188 68960 25194 68972
rect 28258 68960 28264 68972
rect 28316 68960 28322 69012
rect 46566 68960 46572 69012
rect 46624 69000 46630 69012
rect 52822 69000 52828 69012
rect 46624 68972 52828 69000
rect 46624 68960 46630 68972
rect 52822 68960 52828 68972
rect 52880 68960 52886 69012
rect 64138 68960 64144 69012
rect 64196 69000 64202 69012
rect 66990 69000 66996 69012
rect 64196 68972 66996 69000
rect 64196 68960 64202 68972
rect 66990 68960 66996 68972
rect 67048 68960 67054 69012
rect 41874 68892 41880 68944
rect 41932 68932 41938 68944
rect 41932 68904 46980 68932
rect 41932 68892 41938 68904
rect 46477 68867 46535 68873
rect 46477 68833 46489 68867
rect 46523 68864 46535 68867
rect 46750 68864 46756 68876
rect 46523 68836 46756 68864
rect 46523 68833 46535 68836
rect 46477 68827 46535 68833
rect 46750 68824 46756 68836
rect 46808 68824 46814 68876
rect 46952 68873 46980 68904
rect 56686 68892 56692 68944
rect 56744 68932 56750 68944
rect 56744 68904 57100 68932
rect 56744 68892 56750 68904
rect 46937 68867 46995 68873
rect 46937 68833 46949 68867
rect 46983 68833 46995 68867
rect 46937 68827 46995 68833
rect 50985 68867 51043 68873
rect 50985 68833 50997 68867
rect 51031 68864 51043 68867
rect 51258 68864 51264 68876
rect 51031 68836 51264 68864
rect 51031 68833 51043 68836
rect 50985 68827 51043 68833
rect 51258 68824 51264 68836
rect 51316 68824 51322 68876
rect 51534 68864 51540 68876
rect 51495 68836 51540 68864
rect 51534 68824 51540 68836
rect 51592 68824 51598 68876
rect 56229 68867 56287 68873
rect 56229 68833 56241 68867
rect 56275 68864 56287 68867
rect 56962 68864 56968 68876
rect 56275 68836 56968 68864
rect 56275 68833 56287 68836
rect 56229 68827 56287 68833
rect 56962 68824 56968 68836
rect 57020 68824 57026 68876
rect 57072 68873 57100 68904
rect 57057 68867 57115 68873
rect 57057 68833 57069 68867
rect 57103 68833 57115 68867
rect 57057 68827 57115 68833
rect 48777 68799 48835 68805
rect 48777 68765 48789 68799
rect 48823 68796 48835 68799
rect 49142 68796 49148 68808
rect 48823 68768 49148 68796
rect 48823 68765 48835 68768
rect 48777 68759 48835 68765
rect 49142 68756 49148 68768
rect 49200 68756 49206 68808
rect 58894 68796 58900 68808
rect 58855 68768 58900 68796
rect 58894 68756 58900 68768
rect 58952 68756 58958 68808
rect 46661 68731 46719 68737
rect 46661 68697 46673 68731
rect 46707 68697 46719 68731
rect 51166 68728 51172 68740
rect 51127 68700 51172 68728
rect 46661 68691 46719 68697
rect 40678 68620 40684 68672
rect 40736 68660 40742 68672
rect 46566 68660 46572 68672
rect 40736 68632 46572 68660
rect 40736 68620 40742 68632
rect 46566 68620 46572 68632
rect 46624 68620 46630 68672
rect 46676 68660 46704 68691
rect 51166 68688 51172 68700
rect 51224 68688 51230 68740
rect 56410 68728 56416 68740
rect 56371 68700 56416 68728
rect 56410 68688 56416 68700
rect 56468 68688 56474 68740
rect 63126 68728 63132 68740
rect 58912 68700 63132 68728
rect 48869 68663 48927 68669
rect 48869 68660 48881 68663
rect 46676 68632 48881 68660
rect 48869 68629 48881 68632
rect 48915 68629 48927 68663
rect 48869 68623 48927 68629
rect 53282 68620 53288 68672
rect 53340 68660 53346 68672
rect 58912 68660 58940 68700
rect 63126 68688 63132 68700
rect 63184 68688 63190 68740
rect 53340 68632 58940 68660
rect 58989 68663 59047 68669
rect 53340 68620 53346 68632
rect 58989 68629 59001 68663
rect 59035 68660 59047 68663
rect 59170 68660 59176 68672
rect 59035 68632 59176 68660
rect 59035 68629 59047 68632
rect 58989 68623 59047 68629
rect 59170 68620 59176 68632
rect 59228 68620 59234 68672
rect 1104 68570 68816 68592
rect 1104 68518 19574 68570
rect 19626 68518 19638 68570
rect 19690 68518 19702 68570
rect 19754 68518 19766 68570
rect 19818 68518 19830 68570
rect 19882 68518 50294 68570
rect 50346 68518 50358 68570
rect 50410 68518 50422 68570
rect 50474 68518 50486 68570
rect 50538 68518 50550 68570
rect 50602 68518 68816 68570
rect 1104 68496 68816 68518
rect 16758 68416 16764 68468
rect 16816 68456 16822 68468
rect 33134 68456 33140 68468
rect 16816 68428 33140 68456
rect 16816 68416 16822 68428
rect 33134 68416 33140 68428
rect 33192 68416 33198 68468
rect 38562 68416 38568 68468
rect 38620 68456 38626 68468
rect 51166 68456 51172 68468
rect 38620 68428 45554 68456
rect 51127 68428 51172 68456
rect 38620 68416 38626 68428
rect 6454 68348 6460 68400
rect 6512 68388 6518 68400
rect 22738 68388 22744 68400
rect 6512 68360 22744 68388
rect 6512 68348 6518 68360
rect 22738 68348 22744 68360
rect 22796 68348 22802 68400
rect 24118 68348 24124 68400
rect 24176 68388 24182 68400
rect 44450 68388 44456 68400
rect 24176 68360 44456 68388
rect 24176 68348 24182 68360
rect 44450 68348 44456 68360
rect 44508 68348 44514 68400
rect 45526 68388 45554 68428
rect 51166 68416 51172 68428
rect 51224 68416 51230 68468
rect 54110 68456 54116 68468
rect 51276 68428 54116 68456
rect 51276 68388 51304 68428
rect 54110 68416 54116 68428
rect 54168 68416 54174 68468
rect 56410 68456 56416 68468
rect 56371 68428 56416 68456
rect 56410 68416 56416 68428
rect 56468 68416 56474 68468
rect 45526 68360 51304 68388
rect 53374 68348 53380 68400
rect 53432 68388 53438 68400
rect 65334 68388 65340 68400
rect 53432 68360 65340 68388
rect 53432 68348 53438 68360
rect 65334 68348 65340 68360
rect 65392 68348 65398 68400
rect 23198 68280 23204 68332
rect 23256 68320 23262 68332
rect 29638 68320 29644 68332
rect 23256 68292 29644 68320
rect 23256 68280 23262 68292
rect 29638 68280 29644 68292
rect 29696 68280 29702 68332
rect 49142 68280 49148 68332
rect 49200 68320 49206 68332
rect 51077 68323 51135 68329
rect 51077 68320 51089 68323
rect 49200 68292 51089 68320
rect 49200 68280 49206 68292
rect 51077 68289 51089 68292
rect 51123 68320 51135 68323
rect 56321 68323 56379 68329
rect 56321 68320 56333 68323
rect 51123 68292 56333 68320
rect 51123 68289 51135 68292
rect 51077 68283 51135 68289
rect 56321 68289 56333 68292
rect 56367 68289 56379 68323
rect 58986 68320 58992 68332
rect 58947 68292 58992 68320
rect 56321 68283 56379 68289
rect 56336 68252 56364 68283
rect 58986 68280 58992 68292
rect 59044 68280 59050 68332
rect 58894 68252 58900 68264
rect 56336 68224 58900 68252
rect 58894 68212 58900 68224
rect 58952 68212 58958 68264
rect 59170 68252 59176 68264
rect 59131 68224 59176 68252
rect 59170 68212 59176 68224
rect 59228 68212 59234 68264
rect 60829 68255 60887 68261
rect 60829 68221 60841 68255
rect 60875 68252 60887 68255
rect 68278 68252 68284 68264
rect 60875 68224 68284 68252
rect 60875 68221 60887 68224
rect 60829 68215 60887 68221
rect 68278 68212 68284 68224
rect 68336 68212 68342 68264
rect 3878 68076 3884 68128
rect 3936 68116 3942 68128
rect 5534 68116 5540 68128
rect 3936 68088 5540 68116
rect 3936 68076 3942 68088
rect 5534 68076 5540 68088
rect 5592 68076 5598 68128
rect 30282 68076 30288 68128
rect 30340 68116 30346 68128
rect 31110 68116 31116 68128
rect 30340 68088 31116 68116
rect 30340 68076 30346 68088
rect 31110 68076 31116 68088
rect 31168 68076 31174 68128
rect 37918 68076 37924 68128
rect 37976 68116 37982 68128
rect 39298 68116 39304 68128
rect 37976 68088 39304 68116
rect 37976 68076 37982 68088
rect 39298 68076 39304 68088
rect 39356 68076 39362 68128
rect 58618 68076 58624 68128
rect 58676 68116 58682 68128
rect 60550 68116 60556 68128
rect 58676 68088 60556 68116
rect 58676 68076 58682 68088
rect 60550 68076 60556 68088
rect 60608 68076 60614 68128
rect 67726 68076 67732 68128
rect 67784 68116 67790 68128
rect 69198 68116 69204 68128
rect 67784 68088 69204 68116
rect 67784 68076 67790 68088
rect 69198 68076 69204 68088
rect 69256 68076 69262 68128
rect 1104 68026 68816 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 34934 68026
rect 34986 67974 34998 68026
rect 35050 67974 35062 68026
rect 35114 67974 35126 68026
rect 35178 67974 35190 68026
rect 35242 67974 65654 68026
rect 65706 67974 65718 68026
rect 65770 67974 65782 68026
rect 65834 67974 65846 68026
rect 65898 67974 65910 68026
rect 65962 67974 68816 68026
rect 1104 67952 68816 67974
rect 60918 67708 60924 67720
rect 60879 67680 60924 67708
rect 60918 67668 60924 67680
rect 60976 67668 60982 67720
rect 43162 67600 43168 67652
rect 43220 67640 43226 67652
rect 44174 67640 44180 67652
rect 43220 67612 44180 67640
rect 43220 67600 43226 67612
rect 44174 67600 44180 67612
rect 44232 67600 44238 67652
rect 61102 67640 61108 67652
rect 61063 67612 61108 67640
rect 61102 67600 61108 67612
rect 61160 67600 61166 67652
rect 62758 67640 62764 67652
rect 62719 67612 62764 67640
rect 62758 67600 62764 67612
rect 62816 67600 62822 67652
rect 1104 67482 68816 67504
rect 1104 67430 19574 67482
rect 19626 67430 19638 67482
rect 19690 67430 19702 67482
rect 19754 67430 19766 67482
rect 19818 67430 19830 67482
rect 19882 67430 50294 67482
rect 50346 67430 50358 67482
rect 50410 67430 50422 67482
rect 50474 67430 50486 67482
rect 50538 67430 50550 67482
rect 50602 67430 68816 67482
rect 1104 67408 68816 67430
rect 60645 67371 60703 67377
rect 60645 67337 60657 67371
rect 60691 67368 60703 67371
rect 61102 67368 61108 67380
rect 60691 67340 61108 67368
rect 60691 67337 60703 67340
rect 60645 67331 60703 67337
rect 61102 67328 61108 67340
rect 61160 67328 61166 67380
rect 58894 67192 58900 67244
rect 58952 67232 58958 67244
rect 60553 67235 60611 67241
rect 60553 67232 60565 67235
rect 58952 67204 60565 67232
rect 58952 67192 58958 67204
rect 60553 67201 60565 67204
rect 60599 67201 60611 67235
rect 60553 67195 60611 67201
rect 60918 67192 60924 67244
rect 60976 67232 60982 67244
rect 61381 67235 61439 67241
rect 61381 67232 61393 67235
rect 60976 67204 61393 67232
rect 60976 67192 60982 67204
rect 61381 67201 61393 67204
rect 61427 67201 61439 67235
rect 61381 67195 61439 67201
rect 62758 66988 62764 67040
rect 62816 67028 62822 67040
rect 66162 67028 66168 67040
rect 62816 67000 66168 67028
rect 62816 66988 62822 67000
rect 66162 66988 66168 67000
rect 66220 66988 66226 67040
rect 1104 66938 68816 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 68816 66938
rect 1104 66864 68816 66886
rect 37458 66580 37464 66632
rect 37516 66620 37522 66632
rect 37737 66623 37795 66629
rect 37737 66620 37749 66623
rect 37516 66592 37749 66620
rect 37516 66580 37522 66592
rect 37737 66589 37749 66592
rect 37783 66589 37795 66623
rect 37737 66583 37795 66589
rect 43806 66580 43812 66632
rect 43864 66620 43870 66632
rect 44085 66623 44143 66629
rect 44085 66620 44097 66623
rect 43864 66592 44097 66620
rect 43864 66580 43870 66592
rect 44085 66589 44097 66592
rect 44131 66589 44143 66623
rect 44085 66583 44143 66589
rect 1104 66394 68816 66416
rect 1104 66342 19574 66394
rect 19626 66342 19638 66394
rect 19690 66342 19702 66394
rect 19754 66342 19766 66394
rect 19818 66342 19830 66394
rect 19882 66342 50294 66394
rect 50346 66342 50358 66394
rect 50410 66342 50422 66394
rect 50474 66342 50486 66394
rect 50538 66342 50550 66394
rect 50602 66342 68816 66394
rect 1104 66320 68816 66342
rect 37458 66144 37464 66156
rect 37419 66116 37464 66144
rect 37458 66104 37464 66116
rect 37516 66104 37522 66156
rect 43806 66144 43812 66156
rect 43767 66116 43812 66144
rect 43806 66104 43812 66116
rect 43864 66104 43870 66156
rect 37645 66079 37703 66085
rect 37645 66045 37657 66079
rect 37691 66076 37703 66079
rect 37734 66076 37740 66088
rect 37691 66048 37740 66076
rect 37691 66045 37703 66048
rect 37645 66039 37703 66045
rect 37734 66036 37740 66048
rect 37792 66036 37798 66088
rect 38654 66076 38660 66088
rect 38615 66048 38660 66076
rect 38654 66036 38660 66048
rect 38712 66036 38718 66088
rect 43990 66076 43996 66088
rect 43951 66048 43996 66076
rect 43990 66036 43996 66048
rect 44048 66036 44054 66088
rect 45462 66076 45468 66088
rect 45423 66048 45468 66076
rect 45462 66036 45468 66048
rect 45520 66036 45526 66088
rect 1104 65850 68816 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 68816 65850
rect 1104 65776 68816 65798
rect 37734 65736 37740 65748
rect 37695 65708 37740 65736
rect 37734 65696 37740 65708
rect 37792 65696 37798 65748
rect 43809 65739 43867 65745
rect 43809 65705 43821 65739
rect 43855 65736 43867 65739
rect 43990 65736 43996 65748
rect 43855 65708 43996 65736
rect 43855 65705 43867 65708
rect 43809 65699 43867 65705
rect 43990 65696 43996 65708
rect 44048 65696 44054 65748
rect 31386 65560 31392 65612
rect 31444 65600 31450 65612
rect 31444 65572 32352 65600
rect 31444 65560 31450 65572
rect 6730 65492 6736 65544
rect 6788 65532 6794 65544
rect 7009 65535 7067 65541
rect 7009 65532 7021 65535
rect 6788 65504 7021 65532
rect 6788 65492 6794 65504
rect 7009 65501 7021 65504
rect 7055 65501 7067 65535
rect 31846 65532 31852 65544
rect 31807 65504 31852 65532
rect 7009 65495 7067 65501
rect 31846 65492 31852 65504
rect 31904 65492 31910 65544
rect 32324 65541 32352 65572
rect 37660 65572 43760 65600
rect 37660 65541 37688 65572
rect 32309 65535 32367 65541
rect 32309 65501 32321 65535
rect 32355 65501 32367 65535
rect 32309 65495 32367 65501
rect 37645 65535 37703 65541
rect 37645 65501 37657 65535
rect 37691 65501 37703 65535
rect 37645 65495 37703 65501
rect 42610 65492 42616 65544
rect 42668 65532 42674 65544
rect 43732 65541 43760 65572
rect 42889 65535 42947 65541
rect 42889 65532 42901 65535
rect 42668 65504 42901 65532
rect 42668 65492 42674 65504
rect 42889 65501 42901 65504
rect 42935 65501 42947 65535
rect 42889 65495 42947 65501
rect 43717 65535 43775 65541
rect 43717 65501 43729 65535
rect 43763 65532 43775 65535
rect 43898 65532 43904 65544
rect 43763 65504 43904 65532
rect 43763 65501 43775 65504
rect 43717 65495 43775 65501
rect 43898 65492 43904 65504
rect 43956 65492 43962 65544
rect 32585 65467 32643 65473
rect 32585 65433 32597 65467
rect 32631 65464 32643 65467
rect 43530 65464 43536 65476
rect 32631 65436 43536 65464
rect 32631 65433 32643 65436
rect 32585 65427 32643 65433
rect 43530 65424 43536 65436
rect 43588 65424 43594 65476
rect 1104 65306 68816 65328
rect 1104 65254 19574 65306
rect 19626 65254 19638 65306
rect 19690 65254 19702 65306
rect 19754 65254 19766 65306
rect 19818 65254 19830 65306
rect 19882 65254 50294 65306
rect 50346 65254 50358 65306
rect 50410 65254 50422 65306
rect 50474 65254 50486 65306
rect 50538 65254 50550 65306
rect 50602 65254 68816 65306
rect 1104 65232 68816 65254
rect 30926 65084 30932 65136
rect 30984 65124 30990 65136
rect 31481 65127 31539 65133
rect 31481 65124 31493 65127
rect 30984 65096 31493 65124
rect 30984 65084 30990 65096
rect 31481 65093 31493 65096
rect 31527 65124 31539 65127
rect 32309 65127 32367 65133
rect 32309 65124 32321 65127
rect 31527 65096 32321 65124
rect 31527 65093 31539 65096
rect 31481 65087 31539 65093
rect 32309 65093 32321 65096
rect 32355 65093 32367 65127
rect 32309 65087 32367 65093
rect 6730 65056 6736 65068
rect 6691 65028 6736 65056
rect 6730 65016 6736 65028
rect 6788 65016 6794 65068
rect 31386 65056 31392 65068
rect 31347 65028 31392 65056
rect 31386 65016 31392 65028
rect 31444 65016 31450 65068
rect 42610 65056 42616 65068
rect 42571 65028 42616 65056
rect 42610 65016 42616 65028
rect 42668 65016 42674 65068
rect 6914 64948 6920 65000
rect 6972 64988 6978 65000
rect 7193 64991 7251 64997
rect 6972 64960 7017 64988
rect 6972 64948 6978 64960
rect 7193 64957 7205 64991
rect 7239 64957 7251 64991
rect 7193 64951 7251 64957
rect 30929 64991 30987 64997
rect 30929 64957 30941 64991
rect 30975 64988 30987 64991
rect 32125 64991 32183 64997
rect 32125 64988 32137 64991
rect 30975 64960 32137 64988
rect 30975 64957 30987 64960
rect 30929 64951 30987 64957
rect 32125 64957 32137 64960
rect 32171 64957 32183 64991
rect 33134 64988 33140 65000
rect 33095 64960 33140 64988
rect 32125 64951 32183 64957
rect 5534 64880 5540 64932
rect 5592 64920 5598 64932
rect 7208 64920 7236 64951
rect 33134 64948 33140 64960
rect 33192 64948 33198 65000
rect 42794 64988 42800 65000
rect 42755 64960 42800 64988
rect 42794 64948 42800 64960
rect 42852 64948 42858 65000
rect 44174 64988 44180 65000
rect 44135 64960 44180 64988
rect 44174 64948 44180 64960
rect 44232 64948 44238 65000
rect 5592 64892 7236 64920
rect 5592 64880 5598 64892
rect 55950 64852 55956 64864
rect 55911 64824 55956 64852
rect 55950 64812 55956 64824
rect 56008 64812 56014 64864
rect 1104 64762 68816 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 34934 64762
rect 34986 64710 34998 64762
rect 35050 64710 35062 64762
rect 35114 64710 35126 64762
rect 35178 64710 35190 64762
rect 35242 64710 65654 64762
rect 65706 64710 65718 64762
rect 65770 64710 65782 64762
rect 65834 64710 65846 64762
rect 65898 64710 65910 64762
rect 65962 64710 68816 64762
rect 1104 64688 68816 64710
rect 6914 64608 6920 64660
rect 6972 64648 6978 64660
rect 7101 64651 7159 64657
rect 7101 64648 7113 64651
rect 6972 64620 7113 64648
rect 6972 64608 6978 64620
rect 7101 64617 7113 64620
rect 7147 64617 7159 64651
rect 30466 64648 30472 64660
rect 30427 64620 30472 64648
rect 7101 64611 7159 64617
rect 30466 64608 30472 64620
rect 30524 64608 30530 64660
rect 30926 64648 30932 64660
rect 30887 64620 30932 64648
rect 30926 64608 30932 64620
rect 30984 64608 30990 64660
rect 42794 64648 42800 64660
rect 42755 64620 42800 64648
rect 42794 64608 42800 64620
rect 42852 64608 42858 64660
rect 30484 64580 30512 64608
rect 31021 64583 31079 64589
rect 31021 64580 31033 64583
rect 30484 64552 31033 64580
rect 31021 64549 31033 64552
rect 31067 64549 31079 64583
rect 31202 64580 31208 64592
rect 31163 64552 31208 64580
rect 31021 64543 31079 64549
rect 31202 64540 31208 64552
rect 31260 64540 31266 64592
rect 31588 64552 32168 64580
rect 4614 64472 4620 64524
rect 4672 64512 4678 64524
rect 31588 64512 31616 64552
rect 4672 64484 31616 64512
rect 31665 64515 31723 64521
rect 4672 64472 4678 64484
rect 31665 64481 31677 64515
rect 31711 64512 31723 64515
rect 31846 64512 31852 64524
rect 31711 64484 31852 64512
rect 31711 64481 31723 64484
rect 31665 64475 31723 64481
rect 31846 64472 31852 64484
rect 31904 64472 31910 64524
rect 32140 64521 32168 64552
rect 32125 64515 32183 64521
rect 32125 64481 32137 64515
rect 32171 64481 32183 64515
rect 32125 64475 32183 64481
rect 55677 64515 55735 64521
rect 55677 64481 55689 64515
rect 55723 64512 55735 64515
rect 55950 64512 55956 64524
rect 55723 64484 55956 64512
rect 55723 64481 55735 64484
rect 55677 64475 55735 64481
rect 55950 64472 55956 64484
rect 56008 64472 56014 64524
rect 57517 64515 57575 64521
rect 57517 64481 57529 64515
rect 57563 64512 57575 64515
rect 64138 64512 64144 64524
rect 57563 64484 64144 64512
rect 57563 64481 57575 64484
rect 57517 64475 57575 64481
rect 64138 64472 64144 64484
rect 64196 64472 64202 64524
rect 7009 64447 7067 64453
rect 7009 64413 7021 64447
rect 7055 64444 7067 64447
rect 7190 64444 7196 64456
rect 7055 64416 7196 64444
rect 7055 64413 7067 64416
rect 7009 64407 7067 64413
rect 7190 64404 7196 64416
rect 7248 64404 7254 64456
rect 29730 64444 29736 64456
rect 29691 64416 29736 64444
rect 29730 64404 29736 64416
rect 29788 64404 29794 64456
rect 30193 64447 30251 64453
rect 30193 64413 30205 64447
rect 30239 64444 30251 64447
rect 31570 64444 31576 64456
rect 30239 64416 31576 64444
rect 30239 64413 30251 64416
rect 30193 64407 30251 64413
rect 31570 64404 31576 64416
rect 31628 64404 31634 64456
rect 33965 64447 34023 64453
rect 33965 64413 33977 64447
rect 34011 64444 34023 64447
rect 34054 64444 34060 64456
rect 34011 64416 34060 64444
rect 34011 64413 34023 64416
rect 33965 64407 34023 64413
rect 34054 64404 34060 64416
rect 34112 64404 34118 64456
rect 34146 64404 34152 64456
rect 34204 64444 34210 64456
rect 42705 64447 42763 64453
rect 34204 64416 34249 64444
rect 34204 64404 34210 64416
rect 42705 64413 42717 64447
rect 42751 64444 42763 64447
rect 43898 64444 43904 64456
rect 42751 64416 43904 64444
rect 42751 64413 42763 64416
rect 42705 64407 42763 64413
rect 43898 64404 43904 64416
rect 43956 64404 43962 64456
rect 30834 64376 30840 64388
rect 30795 64348 30840 64376
rect 30834 64336 30840 64348
rect 30892 64336 30898 64388
rect 31205 64379 31263 64385
rect 31205 64345 31217 64379
rect 31251 64345 31263 64379
rect 31205 64339 31263 64345
rect 31849 64379 31907 64385
rect 31849 64345 31861 64379
rect 31895 64376 31907 64379
rect 33226 64376 33232 64388
rect 31895 64348 33232 64376
rect 31895 64345 31907 64348
rect 31849 64339 31907 64345
rect 31220 64308 31248 64339
rect 33226 64336 33232 64348
rect 33284 64336 33290 64388
rect 55858 64376 55864 64388
rect 55819 64348 55864 64376
rect 55858 64336 55864 64348
rect 55916 64336 55922 64388
rect 34057 64311 34115 64317
rect 34057 64308 34069 64311
rect 31220 64280 34069 64308
rect 34057 64277 34069 64280
rect 34103 64277 34115 64311
rect 34057 64271 34115 64277
rect 1104 64218 68816 64240
rect 1104 64166 19574 64218
rect 19626 64166 19638 64218
rect 19690 64166 19702 64218
rect 19754 64166 19766 64218
rect 19818 64166 19830 64218
rect 19882 64166 50294 64218
rect 50346 64166 50358 64218
rect 50410 64166 50422 64218
rect 50474 64166 50486 64218
rect 50538 64166 50550 64218
rect 50602 64166 68816 64218
rect 1104 64144 68816 64166
rect 30834 64064 30840 64116
rect 30892 64104 30898 64116
rect 32582 64104 32588 64116
rect 30892 64076 32588 64104
rect 30892 64064 30898 64076
rect 32582 64064 32588 64076
rect 32640 64064 32646 64116
rect 55677 64107 55735 64113
rect 55677 64073 55689 64107
rect 55723 64104 55735 64107
rect 55858 64104 55864 64116
rect 55723 64076 55864 64104
rect 55723 64073 55735 64076
rect 55677 64067 55735 64073
rect 55858 64064 55864 64076
rect 55916 64064 55922 64116
rect 28721 64039 28779 64045
rect 28721 64005 28733 64039
rect 28767 64036 28779 64039
rect 29457 64039 29515 64045
rect 29457 64036 29469 64039
rect 28767 64008 29469 64036
rect 28767 64005 28779 64008
rect 28721 63999 28779 64005
rect 29457 64005 29469 64008
rect 29503 64005 29515 64039
rect 31110 64036 31116 64048
rect 31071 64008 31116 64036
rect 29457 63999 29515 64005
rect 31110 63996 31116 64008
rect 31168 63996 31174 64048
rect 33965 64039 34023 64045
rect 33965 64005 33977 64039
rect 34011 64036 34023 64039
rect 37918 64036 37924 64048
rect 34011 64008 37924 64036
rect 34011 64005 34023 64008
rect 33965 63999 34023 64005
rect 37918 63996 37924 64008
rect 37976 63996 37982 64048
rect 28629 63971 28687 63977
rect 28629 63937 28641 63971
rect 28675 63968 28687 63971
rect 28675 63940 28764 63968
rect 28675 63937 28687 63940
rect 28629 63931 28687 63937
rect 28736 63912 28764 63940
rect 31570 63928 31576 63980
rect 31628 63968 31634 63980
rect 32125 63971 32183 63977
rect 32125 63968 32137 63971
rect 31628 63940 32137 63968
rect 31628 63928 31634 63940
rect 32125 63937 32137 63940
rect 32171 63937 32183 63971
rect 55582 63968 55588 63980
rect 55543 63940 55588 63968
rect 32125 63931 32183 63937
rect 55582 63928 55588 63940
rect 55640 63928 55646 63980
rect 28718 63860 28724 63912
rect 28776 63860 28782 63912
rect 29273 63903 29331 63909
rect 29273 63869 29285 63903
rect 29319 63900 29331 63903
rect 29730 63900 29736 63912
rect 29319 63872 29736 63900
rect 29319 63869 29331 63872
rect 29273 63863 29331 63869
rect 29730 63860 29736 63872
rect 29788 63860 29794 63912
rect 32306 63900 32312 63912
rect 32267 63872 32312 63900
rect 32306 63860 32312 63872
rect 32364 63860 32370 63912
rect 58066 63764 58072 63776
rect 58027 63736 58072 63764
rect 58066 63724 58072 63736
rect 58124 63724 58130 63776
rect 1104 63674 68816 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 34934 63674
rect 34986 63622 34998 63674
rect 35050 63622 35062 63674
rect 35114 63622 35126 63674
rect 35178 63622 35190 63674
rect 35242 63622 65654 63674
rect 65706 63622 65718 63674
rect 65770 63622 65782 63674
rect 65834 63622 65846 63674
rect 65898 63622 65910 63674
rect 65962 63622 68816 63674
rect 1104 63600 68816 63622
rect 28718 63520 28724 63572
rect 28776 63560 28782 63572
rect 30650 63560 30656 63572
rect 28776 63532 30656 63560
rect 28776 63520 28782 63532
rect 30650 63520 30656 63532
rect 30708 63520 30714 63572
rect 33226 63492 33232 63504
rect 33187 63464 33232 63492
rect 33226 63452 33232 63464
rect 33284 63452 33290 63504
rect 29638 63384 29644 63436
rect 29696 63424 29702 63436
rect 31297 63427 31355 63433
rect 31297 63424 31309 63427
rect 29696 63396 31309 63424
rect 29696 63384 29702 63396
rect 31297 63393 31309 63396
rect 31343 63393 31355 63427
rect 31297 63387 31355 63393
rect 57609 63427 57667 63433
rect 57609 63393 57621 63427
rect 57655 63424 57667 63427
rect 58066 63424 58072 63436
rect 57655 63396 58072 63424
rect 57655 63393 57667 63396
rect 57609 63387 57667 63393
rect 58066 63384 58072 63396
rect 58124 63384 58130 63436
rect 59078 63424 59084 63436
rect 59039 63396 59084 63424
rect 59078 63384 59084 63396
rect 59136 63384 59142 63436
rect 30650 63356 30656 63368
rect 30611 63328 30656 63356
rect 30650 63316 30656 63328
rect 30708 63316 30714 63368
rect 31202 63316 31208 63368
rect 31260 63356 31266 63368
rect 31553 63359 31611 63365
rect 31553 63356 31565 63359
rect 31260 63328 31565 63356
rect 31260 63316 31266 63328
rect 31553 63325 31565 63328
rect 31599 63325 31611 63359
rect 33134 63356 33140 63368
rect 33047 63328 33140 63356
rect 31553 63319 31611 63325
rect 33134 63316 33140 63328
rect 33192 63356 33198 63368
rect 44174 63356 44180 63368
rect 33192 63328 44180 63356
rect 33192 63316 33198 63328
rect 44174 63316 44180 63328
rect 44232 63316 44238 63368
rect 49694 63316 49700 63368
rect 49752 63356 49758 63368
rect 50341 63359 50399 63365
rect 50341 63356 50353 63359
rect 49752 63328 50353 63356
rect 49752 63316 49758 63328
rect 50341 63325 50353 63328
rect 50387 63325 50399 63359
rect 50341 63319 50399 63325
rect 30745 63291 30803 63297
rect 30745 63257 30757 63291
rect 30791 63288 30803 63291
rect 32306 63288 32312 63300
rect 30791 63260 32312 63288
rect 30791 63257 30803 63260
rect 30745 63251 30803 63257
rect 32306 63248 32312 63260
rect 32364 63248 32370 63300
rect 57793 63291 57851 63297
rect 57793 63257 57805 63291
rect 57839 63288 57851 63291
rect 57974 63288 57980 63300
rect 57839 63260 57980 63288
rect 57839 63257 57851 63260
rect 57793 63251 57851 63257
rect 57974 63248 57980 63260
rect 58032 63248 58038 63300
rect 32582 63180 32588 63232
rect 32640 63220 32646 63232
rect 32677 63223 32735 63229
rect 32677 63220 32689 63223
rect 32640 63192 32689 63220
rect 32640 63180 32646 63192
rect 32677 63189 32689 63192
rect 32723 63189 32735 63223
rect 32677 63183 32735 63189
rect 1104 63130 68816 63152
rect 1104 63078 19574 63130
rect 19626 63078 19638 63130
rect 19690 63078 19702 63130
rect 19754 63078 19766 63130
rect 19818 63078 19830 63130
rect 19882 63078 50294 63130
rect 50346 63078 50358 63130
rect 50410 63078 50422 63130
rect 50474 63078 50486 63130
rect 50538 63078 50550 63130
rect 50602 63078 68816 63130
rect 1104 63056 68816 63078
rect 49142 63016 49148 63028
rect 49103 62988 49148 63016
rect 49142 62976 49148 62988
rect 49200 62976 49206 63028
rect 57974 63016 57980 63028
rect 57935 62988 57980 63016
rect 57974 62976 57980 62988
rect 58032 62976 58038 63028
rect 48961 62883 49019 62889
rect 48961 62849 48973 62883
rect 49007 62880 49019 62883
rect 49510 62880 49516 62892
rect 49007 62852 49516 62880
rect 49007 62849 49019 62852
rect 48961 62843 49019 62849
rect 49510 62840 49516 62852
rect 49568 62840 49574 62892
rect 49694 62880 49700 62892
rect 49655 62852 49700 62880
rect 49694 62840 49700 62852
rect 49752 62840 49758 62892
rect 57885 62883 57943 62889
rect 57885 62849 57897 62883
rect 57931 62880 57943 62883
rect 64506 62880 64512 62892
rect 57931 62852 64512 62880
rect 57931 62849 57943 62852
rect 57885 62843 57943 62849
rect 64506 62840 64512 62852
rect 64564 62880 64570 62892
rect 64969 62883 65027 62889
rect 64969 62880 64981 62883
rect 64564 62852 64981 62880
rect 64564 62840 64570 62852
rect 64969 62849 64981 62852
rect 65015 62849 65027 62883
rect 64969 62843 65027 62849
rect 31573 62815 31631 62821
rect 31573 62781 31585 62815
rect 31619 62812 31631 62815
rect 32125 62815 32183 62821
rect 32125 62812 32137 62815
rect 31619 62784 32137 62812
rect 31619 62781 31631 62784
rect 31573 62775 31631 62781
rect 32125 62781 32137 62784
rect 32171 62781 32183 62815
rect 32125 62775 32183 62781
rect 32309 62815 32367 62821
rect 32309 62781 32321 62815
rect 32355 62812 32367 62815
rect 32398 62812 32404 62824
rect 32355 62784 32404 62812
rect 32355 62781 32367 62784
rect 32309 62775 32367 62781
rect 32398 62772 32404 62784
rect 32456 62772 32462 62824
rect 32585 62815 32643 62821
rect 32585 62781 32597 62815
rect 32631 62781 32643 62815
rect 32585 62775 32643 62781
rect 49881 62815 49939 62821
rect 49881 62781 49893 62815
rect 49927 62812 49939 62815
rect 50246 62812 50252 62824
rect 49927 62784 50252 62812
rect 49927 62781 49939 62784
rect 49881 62775 49939 62781
rect 30558 62704 30564 62756
rect 30616 62744 30622 62756
rect 32600 62744 32628 62775
rect 50246 62772 50252 62784
rect 50304 62772 50310 62824
rect 50341 62815 50399 62821
rect 50341 62781 50353 62815
rect 50387 62781 50399 62815
rect 50341 62775 50399 62781
rect 30616 62716 32628 62744
rect 30616 62704 30622 62716
rect 49786 62704 49792 62756
rect 49844 62744 49850 62756
rect 50356 62744 50384 62775
rect 49844 62716 50384 62744
rect 49844 62704 49850 62716
rect 65150 62704 65156 62756
rect 65208 62744 65214 62756
rect 65797 62747 65855 62753
rect 65797 62744 65809 62747
rect 65208 62716 65809 62744
rect 65208 62704 65214 62716
rect 65797 62713 65809 62716
rect 65843 62713 65855 62747
rect 65797 62707 65855 62713
rect 46474 62636 46480 62688
rect 46532 62676 46538 62688
rect 46753 62679 46811 62685
rect 46753 62676 46765 62679
rect 46532 62648 46765 62676
rect 46532 62636 46538 62648
rect 46753 62645 46765 62648
rect 46799 62645 46811 62679
rect 46753 62639 46811 62645
rect 65061 62679 65119 62685
rect 65061 62645 65073 62679
rect 65107 62676 65119 62679
rect 65334 62676 65340 62688
rect 65107 62648 65340 62676
rect 65107 62645 65119 62648
rect 65061 62639 65119 62645
rect 65334 62636 65340 62648
rect 65392 62636 65398 62688
rect 1104 62586 68816 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 34934 62586
rect 34986 62534 34998 62586
rect 35050 62534 35062 62586
rect 35114 62534 35126 62586
rect 35178 62534 35190 62586
rect 35242 62534 65654 62586
rect 65706 62534 65718 62586
rect 65770 62534 65782 62586
rect 65834 62534 65846 62586
rect 65898 62534 65910 62586
rect 65962 62534 68816 62586
rect 1104 62512 68816 62534
rect 32398 62472 32404 62484
rect 32359 62444 32404 62472
rect 32398 62432 32404 62444
rect 32456 62432 32462 62484
rect 50246 62472 50252 62484
rect 50207 62444 50252 62472
rect 50246 62432 50252 62444
rect 50304 62432 50310 62484
rect 46474 62336 46480 62348
rect 46435 62308 46480 62336
rect 46474 62296 46480 62308
rect 46532 62296 46538 62348
rect 48222 62336 48228 62348
rect 48183 62308 48228 62336
rect 48222 62296 48228 62308
rect 48280 62296 48286 62348
rect 67450 62336 67456 62348
rect 67411 62308 67456 62336
rect 67450 62296 67456 62308
rect 67508 62296 67514 62348
rect 32309 62271 32367 62277
rect 32309 62237 32321 62271
rect 32355 62268 32367 62271
rect 33134 62268 33140 62280
rect 32355 62240 33140 62268
rect 32355 62237 32367 62240
rect 32309 62231 32367 62237
rect 33134 62228 33140 62240
rect 33192 62228 33198 62280
rect 50157 62271 50215 62277
rect 50157 62237 50169 62271
rect 50203 62237 50215 62271
rect 50157 62231 50215 62237
rect 46658 62200 46664 62212
rect 46619 62172 46664 62200
rect 46658 62160 46664 62172
rect 46716 62160 46722 62212
rect 38470 62092 38476 62144
rect 38528 62132 38534 62144
rect 50172 62132 50200 62231
rect 54478 62228 54484 62280
rect 54536 62268 54542 62280
rect 54665 62271 54723 62277
rect 54665 62268 54677 62271
rect 54536 62240 54677 62268
rect 54536 62228 54542 62240
rect 54665 62237 54677 62240
rect 54711 62237 54723 62271
rect 54665 62231 54723 62237
rect 65061 62271 65119 62277
rect 65061 62237 65073 62271
rect 65107 62268 65119 62271
rect 65613 62271 65671 62277
rect 65613 62268 65625 62271
rect 65107 62240 65625 62268
rect 65107 62237 65119 62240
rect 65061 62231 65119 62237
rect 65613 62237 65625 62240
rect 65659 62237 65671 62271
rect 65613 62231 65671 62237
rect 65794 62200 65800 62212
rect 65755 62172 65800 62200
rect 65794 62160 65800 62172
rect 65852 62160 65858 62212
rect 38528 62104 50200 62132
rect 38528 62092 38534 62104
rect 1104 62042 68816 62064
rect 1104 61990 19574 62042
rect 19626 61990 19638 62042
rect 19690 61990 19702 62042
rect 19754 61990 19766 62042
rect 19818 61990 19830 62042
rect 19882 61990 50294 62042
rect 50346 61990 50358 62042
rect 50410 61990 50422 62042
rect 50474 61990 50486 62042
rect 50538 61990 50550 62042
rect 50602 61990 68816 62042
rect 1104 61968 68816 61990
rect 46658 61928 46664 61940
rect 46619 61900 46664 61928
rect 46658 61888 46664 61900
rect 46716 61888 46722 61940
rect 64601 61931 64659 61937
rect 64601 61897 64613 61931
rect 64647 61928 64659 61931
rect 65794 61928 65800 61940
rect 64647 61900 65800 61928
rect 64647 61897 64659 61900
rect 64601 61891 64659 61897
rect 65794 61888 65800 61900
rect 65852 61888 65858 61940
rect 55582 61860 55588 61872
rect 46584 61832 55588 61860
rect 37274 61752 37280 61804
rect 37332 61792 37338 61804
rect 46584 61801 46612 61832
rect 55582 61820 55588 61832
rect 55640 61820 55646 61872
rect 65334 61860 65340 61872
rect 65295 61832 65340 61860
rect 65334 61820 65340 61832
rect 65392 61820 65398 61872
rect 66993 61863 67051 61869
rect 66993 61829 67005 61863
rect 67039 61860 67051 61863
rect 67726 61860 67732 61872
rect 67039 61832 67732 61860
rect 67039 61829 67051 61832
rect 66993 61823 67051 61829
rect 67726 61820 67732 61832
rect 67784 61820 67790 61872
rect 46569 61795 46627 61801
rect 46569 61792 46581 61795
rect 37332 61764 46581 61792
rect 37332 61752 37338 61764
rect 46569 61761 46581 61764
rect 46615 61761 46627 61795
rect 54478 61792 54484 61804
rect 54439 61764 54484 61792
rect 46569 61755 46627 61761
rect 54478 61752 54484 61764
rect 54536 61752 54542 61804
rect 64506 61792 64512 61804
rect 64467 61764 64512 61792
rect 64506 61752 64512 61764
rect 64564 61752 64570 61804
rect 65150 61792 65156 61804
rect 65111 61764 65156 61792
rect 65150 61752 65156 61764
rect 65208 61752 65214 61804
rect 54662 61724 54668 61736
rect 54623 61696 54668 61724
rect 54662 61684 54668 61696
rect 54720 61684 54726 61736
rect 56321 61727 56379 61733
rect 56321 61693 56333 61727
rect 56367 61724 56379 61727
rect 66070 61724 66076 61736
rect 56367 61696 66076 61724
rect 56367 61693 56379 61696
rect 56321 61687 56379 61693
rect 66070 61684 66076 61696
rect 66128 61684 66134 61736
rect 1104 61498 68816 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 65654 61498
rect 65706 61446 65718 61498
rect 65770 61446 65782 61498
rect 65834 61446 65846 61498
rect 65898 61446 65910 61498
rect 65962 61446 68816 61498
rect 1104 61424 68816 61446
rect 54481 61387 54539 61393
rect 54481 61353 54493 61387
rect 54527 61384 54539 61387
rect 54662 61384 54668 61396
rect 54527 61356 54668 61384
rect 54527 61353 54539 61356
rect 54481 61347 54539 61353
rect 54662 61344 54668 61356
rect 54720 61344 54726 61396
rect 23014 61140 23020 61192
rect 23072 61180 23078 61192
rect 23201 61183 23259 61189
rect 23201 61180 23213 61183
rect 23072 61152 23213 61180
rect 23072 61140 23078 61152
rect 23201 61149 23213 61152
rect 23247 61149 23259 61183
rect 23201 61143 23259 61149
rect 44174 61140 44180 61192
rect 44232 61180 44238 61192
rect 44358 61180 44364 61192
rect 44232 61152 44364 61180
rect 44232 61140 44238 61152
rect 44358 61140 44364 61152
rect 44416 61180 44422 61192
rect 54389 61183 54447 61189
rect 54389 61180 54401 61183
rect 44416 61152 54401 61180
rect 44416 61140 44422 61152
rect 54389 61149 54401 61152
rect 54435 61149 54447 61183
rect 54389 61143 54447 61149
rect 1104 60954 68816 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 68816 60954
rect 1104 60880 68816 60902
rect 23014 60704 23020 60716
rect 22975 60676 23020 60704
rect 23014 60664 23020 60676
rect 23072 60664 23078 60716
rect 1394 60636 1400 60648
rect 1355 60608 1400 60636
rect 1394 60596 1400 60608
rect 1452 60596 1458 60648
rect 1673 60639 1731 60645
rect 1673 60605 1685 60639
rect 1719 60636 1731 60639
rect 23201 60639 23259 60645
rect 1719 60608 6914 60636
rect 1719 60605 1731 60608
rect 1673 60599 1731 60605
rect 6886 60568 6914 60608
rect 23201 60605 23213 60639
rect 23247 60636 23259 60639
rect 23566 60636 23572 60648
rect 23247 60608 23572 60636
rect 23247 60605 23259 60608
rect 23201 60599 23259 60605
rect 23566 60596 23572 60608
rect 23624 60596 23630 60648
rect 23658 60596 23664 60648
rect 23716 60636 23722 60648
rect 23716 60608 23761 60636
rect 23716 60596 23722 60608
rect 34146 60568 34152 60580
rect 6886 60540 34152 60568
rect 34146 60528 34152 60540
rect 34204 60528 34210 60580
rect 22738 60460 22744 60512
rect 22796 60500 22802 60512
rect 23382 60500 23388 60512
rect 22796 60472 23388 60500
rect 22796 60460 22802 60472
rect 23382 60460 23388 60472
rect 23440 60460 23446 60512
rect 1104 60410 68816 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 65654 60410
rect 65706 60358 65718 60410
rect 65770 60358 65782 60410
rect 65834 60358 65846 60410
rect 65898 60358 65910 60410
rect 65962 60358 68816 60410
rect 1104 60336 68816 60358
rect 23566 60296 23572 60308
rect 23527 60268 23572 60296
rect 23566 60256 23572 60268
rect 23624 60256 23630 60308
rect 47210 60188 47216 60240
rect 47268 60228 47274 60240
rect 47268 60200 47624 60228
rect 47268 60188 47274 60200
rect 47596 60169 47624 60200
rect 47581 60163 47639 60169
rect 47581 60129 47593 60163
rect 47627 60129 47639 60163
rect 47581 60123 47639 60129
rect 23477 60095 23535 60101
rect 23477 60061 23489 60095
rect 23523 60092 23535 60095
rect 24854 60092 24860 60104
rect 23523 60064 24860 60092
rect 23523 60061 23535 60064
rect 23477 60055 23535 60061
rect 24854 60052 24860 60064
rect 24912 60052 24918 60104
rect 26970 60092 26976 60104
rect 26931 60064 26976 60092
rect 26970 60052 26976 60064
rect 27028 60052 27034 60104
rect 46661 60095 46719 60101
rect 46661 60061 46673 60095
rect 46707 60092 46719 60095
rect 47121 60095 47179 60101
rect 47121 60092 47133 60095
rect 46707 60064 47133 60092
rect 46707 60061 46719 60064
rect 46661 60055 46719 60061
rect 47121 60061 47133 60064
rect 47167 60061 47179 60095
rect 47121 60055 47179 60061
rect 47305 60027 47363 60033
rect 47305 59993 47317 60027
rect 47351 60024 47363 60027
rect 47670 60024 47676 60036
rect 47351 59996 47676 60024
rect 47351 59993 47363 59996
rect 47305 59987 47363 59993
rect 47670 59984 47676 59996
rect 47728 59984 47734 60036
rect 1104 59866 68816 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 68816 59866
rect 1104 59792 68816 59814
rect 47670 59752 47676 59764
rect 47631 59724 47676 59752
rect 47670 59712 47676 59724
rect 47728 59712 47734 59764
rect 28810 59684 28816 59696
rect 28771 59656 28816 59684
rect 28810 59644 28816 59656
rect 28868 59644 28874 59696
rect 47581 59619 47639 59625
rect 47581 59585 47593 59619
rect 47627 59616 47639 59619
rect 48498 59616 48504 59628
rect 47627 59588 48504 59616
rect 47627 59585 47639 59588
rect 47581 59579 47639 59585
rect 48498 59576 48504 59588
rect 48556 59576 48562 59628
rect 26421 59551 26479 59557
rect 26421 59517 26433 59551
rect 26467 59548 26479 59551
rect 26973 59551 27031 59557
rect 26973 59548 26985 59551
rect 26467 59520 26985 59548
rect 26467 59517 26479 59520
rect 26421 59511 26479 59517
rect 26973 59517 26985 59520
rect 27019 59517 27031 59551
rect 27154 59548 27160 59560
rect 27115 59520 27160 59548
rect 26973 59511 27031 59517
rect 27154 59508 27160 59520
rect 27212 59508 27218 59560
rect 1104 59322 68816 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 65654 59322
rect 65706 59270 65718 59322
rect 65770 59270 65782 59322
rect 65834 59270 65846 59322
rect 65898 59270 65910 59322
rect 65962 59270 68816 59322
rect 1104 59248 68816 59270
rect 26237 59211 26295 59217
rect 26237 59177 26249 59211
rect 26283 59208 26295 59211
rect 27154 59208 27160 59220
rect 26283 59180 27160 59208
rect 26283 59177 26295 59180
rect 26237 59171 26295 59177
rect 27154 59168 27160 59180
rect 27212 59168 27218 59220
rect 26206 59112 27292 59140
rect 26206 59072 26234 59112
rect 6886 59044 26234 59072
rect 26789 59075 26847 59081
rect 3326 58896 3332 58948
rect 3384 58936 3390 58948
rect 6886 58936 6914 59044
rect 26789 59041 26801 59075
rect 26835 59072 26847 59075
rect 26970 59072 26976 59084
rect 26835 59044 26976 59072
rect 26835 59041 26847 59044
rect 26789 59035 26847 59041
rect 26970 59032 26976 59044
rect 27028 59032 27034 59084
rect 27264 59081 27292 59112
rect 27249 59075 27307 59081
rect 27249 59041 27261 59075
rect 27295 59041 27307 59075
rect 27249 59035 27307 59041
rect 24946 58964 24952 59016
rect 25004 59004 25010 59016
rect 26145 59007 26203 59013
rect 26145 59004 26157 59007
rect 25004 58976 26157 59004
rect 25004 58964 25010 58976
rect 26145 58973 26157 58976
rect 26191 58973 26203 59007
rect 26145 58967 26203 58973
rect 3384 58908 6914 58936
rect 26973 58939 27031 58945
rect 3384 58896 3390 58908
rect 26973 58905 26985 58939
rect 27019 58936 27031 58939
rect 27154 58936 27160 58948
rect 27019 58908 27160 58936
rect 27019 58905 27031 58908
rect 26973 58899 27031 58905
rect 27154 58896 27160 58908
rect 27212 58896 27218 58948
rect 1104 58778 68816 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 68816 58778
rect 1104 58704 68816 58726
rect 27154 58664 27160 58676
rect 27115 58636 27160 58664
rect 27154 58624 27160 58636
rect 27212 58624 27218 58676
rect 24854 58488 24860 58540
rect 24912 58528 24918 58540
rect 27065 58531 27123 58537
rect 27065 58528 27077 58531
rect 24912 58500 27077 58528
rect 24912 58488 24918 58500
rect 27065 58497 27077 58500
rect 27111 58528 27123 58531
rect 37918 58528 37924 58540
rect 27111 58500 37924 58528
rect 27111 58497 27123 58500
rect 27065 58491 27123 58497
rect 37918 58488 37924 58500
rect 37976 58528 37982 58540
rect 38470 58528 38476 58540
rect 37976 58500 38476 58528
rect 37976 58488 37982 58500
rect 38470 58488 38476 58500
rect 38528 58488 38534 58540
rect 1104 58234 68816 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 65654 58234
rect 65706 58182 65718 58234
rect 65770 58182 65782 58234
rect 65834 58182 65846 58234
rect 65898 58182 65910 58234
rect 65962 58182 68816 58234
rect 1104 58160 68816 58182
rect 48406 57876 48412 57928
rect 48464 57916 48470 57928
rect 48685 57919 48743 57925
rect 48685 57916 48697 57919
rect 48464 57888 48697 57916
rect 48464 57876 48470 57888
rect 48685 57885 48697 57888
rect 48731 57885 48743 57919
rect 48685 57879 48743 57885
rect 1104 57690 68816 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 68816 57690
rect 1104 57616 68816 57638
rect 48406 57440 48412 57452
rect 48367 57412 48412 57440
rect 48406 57400 48412 57412
rect 48464 57400 48470 57452
rect 48590 57372 48596 57384
rect 48551 57344 48596 57372
rect 48590 57332 48596 57344
rect 48648 57332 48654 57384
rect 48869 57375 48927 57381
rect 48869 57341 48881 57375
rect 48915 57341 48927 57375
rect 48869 57335 48927 57341
rect 48314 57264 48320 57316
rect 48372 57304 48378 57316
rect 48884 57304 48912 57335
rect 48372 57276 48912 57304
rect 48372 57264 48378 57276
rect 1104 57146 68816 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 68816 57146
rect 1104 57072 68816 57094
rect 48590 57032 48596 57044
rect 48551 57004 48596 57032
rect 48590 56992 48596 57004
rect 48648 56992 48654 57044
rect 11054 56856 11060 56908
rect 11112 56896 11118 56908
rect 11609 56899 11667 56905
rect 11609 56896 11621 56899
rect 11112 56868 11621 56896
rect 11112 56856 11118 56868
rect 11609 56865 11621 56868
rect 11655 56865 11667 56899
rect 11609 56859 11667 56865
rect 10689 56831 10747 56837
rect 10689 56797 10701 56831
rect 10735 56828 10747 56831
rect 11149 56831 11207 56837
rect 11149 56828 11161 56831
rect 10735 56800 11161 56828
rect 10735 56797 10747 56800
rect 10689 56791 10747 56797
rect 11149 56797 11161 56800
rect 11195 56797 11207 56831
rect 48498 56828 48504 56840
rect 48411 56800 48504 56828
rect 11149 56791 11207 56797
rect 48498 56788 48504 56800
rect 48556 56828 48562 56840
rect 49050 56828 49056 56840
rect 48556 56800 49056 56828
rect 48556 56788 48562 56800
rect 49050 56788 49056 56800
rect 49108 56788 49114 56840
rect 11330 56760 11336 56772
rect 11291 56732 11336 56760
rect 11330 56720 11336 56732
rect 11388 56720 11394 56772
rect 1104 56602 68816 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 68816 56602
rect 1104 56528 68816 56550
rect 11330 56448 11336 56500
rect 11388 56488 11394 56500
rect 11609 56491 11667 56497
rect 11609 56488 11621 56491
rect 11388 56460 11621 56488
rect 11388 56448 11394 56460
rect 11609 56457 11621 56460
rect 11655 56457 11667 56491
rect 11609 56451 11667 56457
rect 20622 56448 20628 56500
rect 20680 56488 20686 56500
rect 24946 56488 24952 56500
rect 20680 56460 24952 56488
rect 20680 56448 20686 56460
rect 24946 56448 24952 56460
rect 25004 56448 25010 56500
rect 11514 56352 11520 56364
rect 11427 56324 11520 56352
rect 11514 56312 11520 56324
rect 11572 56352 11578 56364
rect 20622 56352 20628 56364
rect 11572 56324 20628 56352
rect 11572 56312 11578 56324
rect 20622 56312 20628 56324
rect 20680 56312 20686 56364
rect 1104 56058 68816 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 68816 56058
rect 1104 55984 68816 56006
rect 57333 55743 57391 55749
rect 57333 55709 57345 55743
rect 57379 55740 57391 55743
rect 57882 55740 57888 55752
rect 57379 55712 57888 55740
rect 57379 55709 57391 55712
rect 57333 55703 57391 55709
rect 57882 55700 57888 55712
rect 57940 55700 57946 55752
rect 2958 55564 2964 55616
rect 3016 55604 3022 55616
rect 33042 55604 33048 55616
rect 3016 55576 33048 55604
rect 3016 55564 3022 55576
rect 33042 55564 33048 55576
rect 33100 55564 33106 55616
rect 1104 55514 68816 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 68816 55514
rect 1104 55440 68816 55462
rect 32769 55335 32827 55341
rect 32769 55301 32781 55335
rect 32815 55332 32827 55335
rect 37369 55335 37427 55341
rect 37369 55332 37381 55335
rect 32815 55304 37381 55332
rect 32815 55301 32827 55304
rect 32769 55295 32827 55301
rect 37369 55301 37381 55304
rect 37415 55301 37427 55335
rect 37369 55295 37427 55301
rect 57057 55335 57115 55341
rect 57057 55301 57069 55335
rect 57103 55332 57115 55335
rect 58069 55335 58127 55341
rect 58069 55332 58081 55335
rect 57103 55304 58081 55332
rect 57103 55301 57115 55304
rect 57057 55295 57115 55301
rect 58069 55301 58081 55304
rect 58115 55301 58127 55335
rect 58069 55295 58127 55301
rect 32582 55264 32588 55276
rect 32543 55236 32588 55264
rect 32582 55224 32588 55236
rect 32640 55224 32646 55276
rect 37274 55264 37280 55276
rect 37235 55236 37280 55264
rect 37274 55224 37280 55236
rect 37332 55224 37338 55276
rect 49050 55224 49056 55276
rect 49108 55264 49114 55276
rect 56965 55267 57023 55273
rect 56965 55264 56977 55267
rect 49108 55236 56977 55264
rect 49108 55224 49114 55236
rect 56965 55233 56977 55236
rect 57011 55233 57023 55267
rect 57882 55264 57888 55276
rect 57843 55236 57888 55264
rect 56965 55227 57023 55233
rect 57882 55224 57888 55236
rect 57940 55224 57946 55276
rect 59725 55267 59783 55273
rect 59725 55233 59737 55267
rect 59771 55264 59783 55267
rect 59771 55236 62068 55264
rect 59771 55233 59783 55236
rect 59725 55227 59783 55233
rect 33042 55196 33048 55208
rect 33003 55168 33048 55196
rect 33042 55156 33048 55168
rect 33100 55156 33106 55208
rect 62040 55196 62068 55236
rect 66070 55196 66076 55208
rect 62040 55168 66076 55196
rect 66070 55156 66076 55168
rect 66128 55156 66134 55208
rect 1104 54970 68816 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 68816 54970
rect 1104 54896 68816 54918
rect 1104 54426 68816 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 68816 54426
rect 1104 54352 68816 54374
rect 2774 54000 2780 54052
rect 2832 54040 2838 54052
rect 5718 54040 5724 54052
rect 2832 54012 5724 54040
rect 2832 54000 2838 54012
rect 5718 54000 5724 54012
rect 5776 54000 5782 54052
rect 27522 53972 27528 53984
rect 27483 53944 27528 53972
rect 27522 53932 27528 53944
rect 27580 53932 27586 53984
rect 38838 53932 38844 53984
rect 38896 53972 38902 53984
rect 39025 53975 39083 53981
rect 39025 53972 39037 53975
rect 38896 53944 39037 53972
rect 38896 53932 38902 53944
rect 39025 53941 39037 53944
rect 39071 53941 39083 53975
rect 51442 53972 51448 53984
rect 51403 53944 51448 53972
rect 39025 53935 39083 53941
rect 51442 53932 51448 53944
rect 51500 53932 51506 53984
rect 66254 53932 66260 53984
rect 66312 53972 66318 53984
rect 67637 53975 67695 53981
rect 67637 53972 67649 53975
rect 66312 53944 67649 53972
rect 66312 53932 66318 53944
rect 67637 53941 67649 53944
rect 67683 53941 67695 53975
rect 67637 53935 67695 53941
rect 1104 53882 68816 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 68816 53882
rect 1104 53808 68816 53830
rect 26206 53672 27660 53700
rect 3510 53592 3516 53644
rect 3568 53632 3574 53644
rect 26206 53632 26234 53672
rect 3568 53604 26234 53632
rect 27157 53635 27215 53641
rect 3568 53592 3574 53604
rect 27157 53601 27169 53635
rect 27203 53632 27215 53635
rect 27522 53632 27528 53644
rect 27203 53604 27528 53632
rect 27203 53601 27215 53604
rect 27157 53595 27215 53601
rect 27522 53592 27528 53604
rect 27580 53592 27586 53644
rect 27632 53641 27660 53672
rect 66162 53660 66168 53712
rect 66220 53700 66226 53712
rect 66220 53672 66760 53700
rect 66220 53660 66226 53672
rect 27617 53635 27675 53641
rect 27617 53601 27629 53635
rect 27663 53601 27675 53635
rect 27617 53595 27675 53601
rect 51169 53635 51227 53641
rect 51169 53601 51181 53635
rect 51215 53632 51227 53635
rect 51442 53632 51448 53644
rect 51215 53604 51448 53632
rect 51215 53601 51227 53604
rect 51169 53595 51227 53601
rect 51442 53592 51448 53604
rect 51500 53592 51506 53644
rect 66254 53632 66260 53644
rect 66215 53604 66260 53632
rect 66254 53592 66260 53604
rect 66312 53592 66318 53644
rect 66732 53641 66760 53672
rect 66717 53635 66775 53641
rect 66717 53601 66729 53635
rect 66763 53601 66775 53635
rect 66717 53595 66775 53601
rect 27341 53499 27399 53505
rect 27341 53465 27353 53499
rect 27387 53496 27399 53499
rect 27890 53496 27896 53508
rect 27387 53468 27896 53496
rect 27387 53465 27399 53468
rect 27341 53459 27399 53465
rect 27890 53456 27896 53468
rect 27948 53456 27954 53508
rect 51350 53496 51356 53508
rect 51311 53468 51356 53496
rect 51350 53456 51356 53468
rect 51408 53456 51414 53508
rect 53009 53499 53067 53505
rect 53009 53465 53021 53499
rect 53055 53496 53067 53499
rect 58618 53496 58624 53508
rect 53055 53468 58624 53496
rect 53055 53465 53067 53468
rect 53009 53459 53067 53465
rect 58618 53456 58624 53468
rect 58676 53456 58682 53508
rect 66438 53496 66444 53508
rect 66399 53468 66444 53496
rect 66438 53456 66444 53468
rect 66496 53456 66502 53508
rect 1104 53338 68816 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 68816 53338
rect 1104 53264 68816 53286
rect 27890 53224 27896 53236
rect 27851 53196 27896 53224
rect 27890 53184 27896 53196
rect 27948 53184 27954 53236
rect 51169 53227 51227 53233
rect 51169 53193 51181 53227
rect 51215 53224 51227 53227
rect 51350 53224 51356 53236
rect 51215 53196 51356 53224
rect 51215 53193 51227 53196
rect 51169 53187 51227 53193
rect 51350 53184 51356 53196
rect 51408 53184 51414 53236
rect 66438 53184 66444 53236
rect 66496 53224 66502 53236
rect 67545 53227 67603 53233
rect 67545 53224 67557 53227
rect 66496 53196 67557 53224
rect 66496 53184 66502 53196
rect 67545 53193 67557 53196
rect 67591 53193 67603 53227
rect 67545 53187 67603 53193
rect 38289 53159 38347 53165
rect 38289 53125 38301 53159
rect 38335 53156 38347 53159
rect 39025 53159 39083 53165
rect 39025 53156 39037 53159
rect 38335 53128 39037 53156
rect 38335 53125 38347 53128
rect 38289 53119 38347 53125
rect 39025 53125 39037 53128
rect 39071 53125 39083 53159
rect 40678 53156 40684 53168
rect 40639 53128 40684 53156
rect 39025 53119 39083 53125
rect 40678 53116 40684 53128
rect 40736 53116 40742 53168
rect 27801 53091 27859 53097
rect 27801 53057 27813 53091
rect 27847 53088 27859 53091
rect 38194 53088 38200 53100
rect 27847 53060 35894 53088
rect 38155 53060 38200 53088
rect 27847 53057 27859 53060
rect 27801 53051 27859 53057
rect 35866 52952 35894 53060
rect 38194 53048 38200 53060
rect 38252 53048 38258 53100
rect 38838 53088 38844 53100
rect 38799 53060 38844 53088
rect 38838 53048 38844 53060
rect 38896 53048 38902 53100
rect 51074 53088 51080 53100
rect 51035 53060 51080 53088
rect 51074 53048 51080 53060
rect 51132 53048 51138 53100
rect 67450 53088 67456 53100
rect 67411 53060 67456 53088
rect 67450 53048 67456 53060
rect 67508 53048 67514 53100
rect 45370 52952 45376 52964
rect 35866 52924 45376 52952
rect 45370 52912 45376 52924
rect 45428 52912 45434 52964
rect 5258 52844 5264 52896
rect 5316 52884 5322 52896
rect 5537 52887 5595 52893
rect 5537 52884 5549 52887
rect 5316 52856 5549 52884
rect 5316 52844 5322 52856
rect 5537 52853 5549 52856
rect 5583 52853 5595 52887
rect 5537 52847 5595 52853
rect 7558 52844 7564 52896
rect 7616 52884 7622 52896
rect 7837 52887 7895 52893
rect 7837 52884 7849 52887
rect 7616 52856 7849 52884
rect 7616 52844 7622 52856
rect 7837 52853 7849 52856
rect 7883 52853 7895 52887
rect 7837 52847 7895 52853
rect 1104 52794 68816 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 68816 52794
rect 1104 52720 68816 52742
rect 5258 52544 5264 52556
rect 5219 52516 5264 52544
rect 5258 52504 5264 52516
rect 5316 52504 5322 52556
rect 5445 52547 5503 52553
rect 5445 52513 5457 52547
rect 5491 52544 5503 52547
rect 5626 52544 5632 52556
rect 5491 52516 5632 52544
rect 5491 52513 5503 52516
rect 5445 52507 5503 52513
rect 5626 52504 5632 52516
rect 5684 52504 5690 52556
rect 5718 52504 5724 52556
rect 5776 52544 5782 52556
rect 5776 52516 5821 52544
rect 5776 52504 5782 52516
rect 8113 52479 8171 52485
rect 8113 52445 8125 52479
rect 8159 52476 8171 52479
rect 11514 52476 11520 52488
rect 8159 52448 11520 52476
rect 8159 52445 8171 52448
rect 8113 52439 8171 52445
rect 11514 52436 11520 52448
rect 11572 52436 11578 52488
rect 7742 52300 7748 52352
rect 7800 52340 7806 52352
rect 8205 52343 8263 52349
rect 8205 52340 8217 52343
rect 7800 52312 8217 52340
rect 7800 52300 7806 52312
rect 8205 52309 8217 52312
rect 8251 52309 8263 52343
rect 8205 52303 8263 52309
rect 1104 52250 68816 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 68816 52250
rect 1104 52176 68816 52198
rect 5626 52096 5632 52148
rect 5684 52136 5690 52148
rect 5721 52139 5779 52145
rect 5721 52136 5733 52139
rect 5684 52108 5733 52136
rect 5684 52096 5690 52108
rect 5721 52105 5733 52108
rect 5767 52105 5779 52139
rect 5721 52099 5779 52105
rect 2958 52028 2964 52080
rect 3016 52068 3022 52080
rect 7742 52068 7748 52080
rect 3016 52040 6914 52068
rect 7703 52040 7748 52068
rect 3016 52028 3022 52040
rect 5629 52003 5687 52009
rect 5629 51969 5641 52003
rect 5675 51969 5687 52003
rect 5629 51963 5687 51969
rect 5644 51864 5672 51963
rect 6886 51932 6914 52040
rect 7742 52028 7748 52040
rect 7800 52028 7806 52080
rect 7558 52000 7564 52012
rect 7519 51972 7564 52000
rect 7558 51960 7564 51972
rect 7616 51960 7622 52012
rect 8021 51935 8079 51941
rect 8021 51932 8033 51935
rect 6886 51904 8033 51932
rect 8021 51901 8033 51904
rect 8067 51901 8079 51935
rect 8021 51895 8079 51901
rect 20898 51864 20904 51876
rect 5644 51836 20904 51864
rect 20898 51824 20904 51836
rect 20956 51824 20962 51876
rect 51350 51756 51356 51808
rect 51408 51796 51414 51808
rect 51629 51799 51687 51805
rect 51629 51796 51641 51799
rect 51408 51768 51641 51796
rect 51408 51756 51414 51768
rect 51629 51765 51641 51768
rect 51675 51765 51687 51799
rect 51629 51759 51687 51765
rect 1104 51706 68816 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 68816 51706
rect 1104 51632 68816 51654
rect 51350 51456 51356 51468
rect 51311 51428 51356 51456
rect 51350 51416 51356 51428
rect 51408 51416 51414 51468
rect 53193 51459 53251 51465
rect 53193 51425 53205 51459
rect 53239 51456 53251 51459
rect 53282 51456 53288 51468
rect 53239 51428 53288 51456
rect 53239 51425 53251 51428
rect 53193 51419 53251 51425
rect 53282 51416 53288 51428
rect 53340 51416 53346 51468
rect 34882 51348 34888 51400
rect 34940 51388 34946 51400
rect 35529 51391 35587 51397
rect 35529 51388 35541 51391
rect 34940 51360 35541 51388
rect 34940 51348 34946 51360
rect 35529 51357 35541 51360
rect 35575 51357 35587 51391
rect 35529 51351 35587 51357
rect 45554 51348 45560 51400
rect 45612 51388 45618 51400
rect 45612 51360 45657 51388
rect 45612 51348 45618 51360
rect 51534 51320 51540 51332
rect 51495 51292 51540 51320
rect 51534 51280 51540 51292
rect 51592 51280 51598 51332
rect 36722 51212 36728 51264
rect 36780 51252 36786 51264
rect 66070 51252 66076 51264
rect 36780 51224 66076 51252
rect 36780 51212 36786 51224
rect 66070 51212 66076 51224
rect 66128 51212 66134 51264
rect 1104 51162 68816 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 68816 51162
rect 1104 51088 68816 51110
rect 51353 51051 51411 51057
rect 51353 51017 51365 51051
rect 51399 51048 51411 51051
rect 51534 51048 51540 51060
rect 51399 51020 51540 51048
rect 51399 51017 51411 51020
rect 51353 51011 51411 51017
rect 51534 51008 51540 51020
rect 51592 51008 51598 51060
rect 3326 50940 3332 50992
rect 3384 50980 3390 50992
rect 36722 50980 36728 50992
rect 3384 50952 36400 50980
rect 36683 50952 36728 50980
rect 3384 50940 3390 50952
rect 34882 50912 34888 50924
rect 34843 50884 34888 50912
rect 34882 50872 34888 50884
rect 34940 50872 34946 50924
rect 35069 50847 35127 50853
rect 35069 50813 35081 50847
rect 35115 50844 35127 50847
rect 35342 50844 35348 50856
rect 35115 50816 35348 50844
rect 35115 50813 35127 50816
rect 35069 50807 35127 50813
rect 35342 50804 35348 50816
rect 35400 50804 35406 50856
rect 36372 50776 36400 50952
rect 36722 50940 36728 50952
rect 36780 50940 36786 50992
rect 45554 50980 45560 50992
rect 45204 50952 45560 50980
rect 45204 50921 45232 50952
rect 45554 50940 45560 50952
rect 45612 50940 45618 50992
rect 45189 50915 45247 50921
rect 45189 50881 45201 50915
rect 45235 50881 45247 50915
rect 45189 50875 45247 50881
rect 51261 50915 51319 50921
rect 51261 50881 51273 50915
rect 51307 50912 51319 50915
rect 53190 50912 53196 50924
rect 51307 50884 53196 50912
rect 51307 50881 51319 50884
rect 51261 50875 51319 50881
rect 53190 50872 53196 50884
rect 53248 50872 53254 50924
rect 45373 50847 45431 50853
rect 45373 50813 45385 50847
rect 45419 50844 45431 50847
rect 45554 50844 45560 50856
rect 45419 50816 45560 50844
rect 45419 50813 45431 50816
rect 45373 50807 45431 50813
rect 45554 50804 45560 50816
rect 45612 50804 45618 50856
rect 45649 50847 45707 50853
rect 45649 50813 45661 50847
rect 45695 50813 45707 50847
rect 45649 50807 45707 50813
rect 45664 50776 45692 50807
rect 36372 50748 45692 50776
rect 63218 50668 63224 50720
rect 63276 50708 63282 50720
rect 63681 50711 63739 50717
rect 63681 50708 63693 50711
rect 63276 50680 63693 50708
rect 63276 50668 63282 50680
rect 63681 50677 63693 50680
rect 63727 50677 63739 50711
rect 63681 50671 63739 50677
rect 1104 50618 68816 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 68816 50618
rect 1104 50544 68816 50566
rect 35342 50504 35348 50516
rect 35303 50476 35348 50504
rect 35342 50464 35348 50476
rect 35400 50464 35406 50516
rect 45554 50464 45560 50516
rect 45612 50504 45618 50516
rect 46017 50507 46075 50513
rect 46017 50504 46029 50507
rect 45612 50476 46029 50504
rect 45612 50464 45618 50476
rect 46017 50473 46029 50476
rect 46063 50473 46075 50507
rect 46017 50467 46075 50473
rect 63218 50368 63224 50380
rect 63179 50340 63224 50368
rect 63218 50328 63224 50340
rect 63276 50328 63282 50380
rect 64782 50368 64788 50380
rect 64743 50340 64788 50368
rect 64782 50328 64788 50340
rect 64840 50328 64846 50380
rect 6914 50260 6920 50312
rect 6972 50300 6978 50312
rect 7193 50303 7251 50309
rect 7193 50300 7205 50303
rect 6972 50272 7205 50300
rect 6972 50260 6978 50272
rect 7193 50269 7205 50272
rect 7239 50269 7251 50303
rect 7193 50263 7251 50269
rect 27430 50260 27436 50312
rect 27488 50300 27494 50312
rect 28721 50303 28779 50309
rect 28721 50300 28733 50303
rect 27488 50272 28733 50300
rect 27488 50260 27494 50272
rect 28721 50269 28733 50272
rect 28767 50269 28779 50303
rect 28721 50263 28779 50269
rect 29730 50260 29736 50312
rect 29788 50300 29794 50312
rect 30285 50303 30343 50309
rect 30285 50300 30297 50303
rect 29788 50272 30297 50300
rect 29788 50260 29794 50272
rect 30285 50269 30297 50272
rect 30331 50269 30343 50303
rect 30285 50263 30343 50269
rect 35253 50303 35311 50309
rect 35253 50269 35265 50303
rect 35299 50300 35311 50303
rect 35434 50300 35440 50312
rect 35299 50272 35440 50300
rect 35299 50269 35311 50272
rect 35253 50263 35311 50269
rect 35434 50260 35440 50272
rect 35492 50300 35498 50312
rect 38194 50300 38200 50312
rect 35492 50272 38200 50300
rect 35492 50260 35498 50272
rect 38194 50260 38200 50272
rect 38252 50260 38258 50312
rect 45925 50303 45983 50309
rect 45925 50269 45937 50303
rect 45971 50300 45983 50303
rect 47578 50300 47584 50312
rect 45971 50272 47584 50300
rect 45971 50269 45983 50272
rect 45925 50263 45983 50269
rect 47578 50260 47584 50272
rect 47636 50260 47642 50312
rect 63402 50232 63408 50244
rect 63363 50204 63408 50232
rect 63402 50192 63408 50204
rect 63460 50192 63466 50244
rect 1104 50074 68816 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 68816 50074
rect 1104 50000 68816 50022
rect 28258 49920 28264 49972
rect 28316 49960 28322 49972
rect 63221 49963 63279 49969
rect 28316 49932 30788 49960
rect 28316 49920 28322 49932
rect 29270 49892 29276 49904
rect 29231 49864 29276 49892
rect 29270 49852 29276 49864
rect 29328 49852 29334 49904
rect 30760 49892 30788 49932
rect 63221 49929 63233 49963
rect 63267 49960 63279 49963
rect 63402 49960 63408 49972
rect 63267 49932 63408 49960
rect 63267 49929 63279 49932
rect 63221 49923 63279 49929
rect 63402 49920 63408 49932
rect 63460 49920 63466 49972
rect 30760 49864 31156 49892
rect 6914 49824 6920 49836
rect 6875 49796 6920 49824
rect 6914 49784 6920 49796
rect 6972 49784 6978 49836
rect 27430 49824 27436 49836
rect 27391 49796 27436 49824
rect 27430 49784 27436 49796
rect 27488 49784 27494 49836
rect 29730 49824 29736 49836
rect 29691 49796 29736 49824
rect 29730 49784 29736 49796
rect 29788 49784 29794 49836
rect 4062 49716 4068 49768
rect 4120 49756 4126 49768
rect 7098 49756 7104 49768
rect 4120 49728 6960 49756
rect 7059 49728 7104 49756
rect 4120 49716 4126 49728
rect 6932 49688 6960 49728
rect 7098 49716 7104 49728
rect 7156 49716 7162 49768
rect 7377 49759 7435 49765
rect 7377 49756 7389 49759
rect 7208 49728 7389 49756
rect 7208 49688 7236 49728
rect 7377 49725 7389 49728
rect 7423 49725 7435 49759
rect 27614 49756 27620 49768
rect 27575 49728 27620 49756
rect 7377 49719 7435 49725
rect 27614 49716 27620 49728
rect 27672 49716 27678 49768
rect 29917 49759 29975 49765
rect 29917 49725 29929 49759
rect 29963 49756 29975 49759
rect 30374 49756 30380 49768
rect 29963 49728 30380 49756
rect 29963 49725 29975 49728
rect 29917 49719 29975 49725
rect 30374 49716 30380 49728
rect 30432 49716 30438 49768
rect 31128 49765 31156 49864
rect 62942 49784 62948 49836
rect 63000 49824 63006 49836
rect 63129 49827 63187 49833
rect 63129 49824 63141 49827
rect 63000 49796 63141 49824
rect 63000 49784 63006 49796
rect 63129 49793 63141 49796
rect 63175 49793 63187 49827
rect 63129 49787 63187 49793
rect 31113 49759 31171 49765
rect 31113 49725 31125 49759
rect 31159 49725 31171 49759
rect 31113 49719 31171 49725
rect 6932 49660 7236 49688
rect 1104 49530 68816 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 68816 49530
rect 1104 49456 68816 49478
rect 7098 49376 7104 49428
rect 7156 49416 7162 49428
rect 7285 49419 7343 49425
rect 7285 49416 7297 49419
rect 7156 49388 7297 49416
rect 7156 49376 7162 49388
rect 7285 49385 7297 49388
rect 7331 49385 7343 49419
rect 7285 49379 7343 49385
rect 27614 49376 27620 49428
rect 27672 49416 27678 49428
rect 28629 49419 28687 49425
rect 28629 49416 28641 49419
rect 27672 49388 28641 49416
rect 27672 49376 27678 49388
rect 28629 49385 28641 49388
rect 28675 49385 28687 49419
rect 30374 49416 30380 49428
rect 30335 49388 30380 49416
rect 28629 49379 28687 49385
rect 30374 49376 30380 49388
rect 30432 49376 30438 49428
rect 7190 49212 7196 49224
rect 7151 49184 7196 49212
rect 7190 49172 7196 49184
rect 7248 49172 7254 49224
rect 28534 49212 28540 49224
rect 28495 49184 28540 49212
rect 28534 49172 28540 49184
rect 28592 49172 28598 49224
rect 30285 49215 30343 49221
rect 30285 49181 30297 49215
rect 30331 49212 30343 49215
rect 41598 49212 41604 49224
rect 30331 49184 41604 49212
rect 30331 49181 30343 49184
rect 30285 49175 30343 49181
rect 41598 49172 41604 49184
rect 41656 49172 41662 49224
rect 53834 49172 53840 49224
rect 53892 49212 53898 49224
rect 54113 49215 54171 49221
rect 54113 49212 54125 49215
rect 53892 49184 54125 49212
rect 53892 49172 53898 49184
rect 54113 49181 54125 49184
rect 54159 49181 54171 49215
rect 54113 49175 54171 49181
rect 1104 48986 68816 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 68816 48986
rect 1104 48912 68816 48934
rect 44358 48764 44364 48816
rect 44416 48804 44422 48816
rect 44453 48807 44511 48813
rect 44453 48804 44465 48807
rect 44416 48776 44465 48804
rect 44416 48764 44422 48776
rect 44453 48773 44465 48776
rect 44499 48773 44511 48807
rect 44453 48767 44511 48773
rect 53285 48807 53343 48813
rect 53285 48773 53297 48807
rect 53331 48804 53343 48807
rect 54021 48807 54079 48813
rect 54021 48804 54033 48807
rect 53331 48776 54033 48804
rect 53331 48773 53343 48776
rect 53285 48767 53343 48773
rect 54021 48773 54033 48776
rect 54067 48773 54079 48807
rect 54021 48767 54079 48773
rect 55677 48807 55735 48813
rect 55677 48773 55689 48807
rect 55723 48804 55735 48807
rect 64690 48804 64696 48816
rect 55723 48776 64696 48804
rect 55723 48773 55735 48776
rect 55677 48767 55735 48773
rect 64690 48764 64696 48776
rect 64748 48764 64754 48816
rect 43533 48739 43591 48745
rect 43533 48705 43545 48739
rect 43579 48705 43591 48739
rect 44174 48736 44180 48748
rect 44135 48708 44180 48736
rect 43533 48699 43591 48705
rect 43548 48668 43576 48699
rect 44174 48696 44180 48708
rect 44232 48736 44238 48748
rect 45189 48739 45247 48745
rect 45189 48736 45201 48739
rect 44232 48708 45201 48736
rect 44232 48696 44238 48708
rect 45189 48705 45201 48708
rect 45235 48705 45247 48739
rect 53190 48736 53196 48748
rect 53151 48708 53196 48736
rect 45189 48699 45247 48705
rect 53190 48696 53196 48708
rect 53248 48696 53254 48748
rect 53834 48736 53840 48748
rect 53795 48708 53840 48736
rect 53834 48696 53840 48708
rect 53892 48696 53898 48748
rect 45465 48671 45523 48677
rect 45465 48668 45477 48671
rect 43548 48640 45477 48668
rect 45465 48637 45477 48640
rect 45511 48637 45523 48671
rect 45465 48631 45523 48637
rect 45480 48600 45508 48631
rect 64506 48600 64512 48612
rect 45480 48572 64512 48600
rect 64506 48560 64512 48572
rect 64564 48600 64570 48612
rect 64690 48600 64696 48612
rect 64564 48572 64696 48600
rect 64564 48560 64570 48572
rect 64690 48560 64696 48572
rect 64748 48560 64754 48612
rect 43622 48532 43628 48544
rect 43583 48504 43628 48532
rect 43622 48492 43628 48504
rect 43680 48492 43686 48544
rect 1104 48442 68816 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 68816 48442
rect 1104 48368 68816 48390
rect 43898 48220 43904 48272
rect 43956 48260 43962 48272
rect 43993 48263 44051 48269
rect 43993 48260 44005 48263
rect 43956 48232 44005 48260
rect 43956 48220 43962 48232
rect 43993 48229 44005 48232
rect 44039 48229 44051 48263
rect 43993 48223 44051 48229
rect 43257 48127 43315 48133
rect 43257 48093 43269 48127
rect 43303 48124 43315 48127
rect 43438 48124 43444 48136
rect 43303 48096 43444 48124
rect 43303 48093 43315 48096
rect 43257 48087 43315 48093
rect 43438 48084 43444 48096
rect 43496 48084 43502 48136
rect 45005 48127 45063 48133
rect 45005 48093 45017 48127
rect 45051 48093 45063 48127
rect 45005 48087 45063 48093
rect 43809 48059 43867 48065
rect 43809 48025 43821 48059
rect 43855 48056 43867 48059
rect 44174 48056 44180 48068
rect 43855 48028 44180 48056
rect 43855 48025 43867 48028
rect 43809 48019 43867 48025
rect 44174 48016 44180 48028
rect 44232 48056 44238 48068
rect 45020 48056 45048 48087
rect 45278 48056 45284 48068
rect 44232 48028 45048 48056
rect 45191 48028 45284 48056
rect 44232 48016 44238 48028
rect 45278 48016 45284 48028
rect 45336 48056 45342 48068
rect 53190 48056 53196 48068
rect 45336 48028 53196 48056
rect 45336 48016 45342 48028
rect 53190 48016 53196 48028
rect 53248 48016 53254 48068
rect 1104 47898 68816 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 68816 47898
rect 1104 47824 68816 47846
rect 43622 47716 43628 47728
rect 43583 47688 43628 47716
rect 43622 47676 43628 47688
rect 43680 47676 43686 47728
rect 64785 47719 64843 47725
rect 64785 47685 64797 47719
rect 64831 47716 64843 47719
rect 65521 47719 65579 47725
rect 65521 47716 65533 47719
rect 64831 47688 65533 47716
rect 64831 47685 64843 47688
rect 64785 47679 64843 47685
rect 65521 47685 65533 47688
rect 65567 47685 65579 47719
rect 65521 47679 65579 47685
rect 43438 47648 43444 47660
rect 43399 47620 43444 47648
rect 43438 47608 43444 47620
rect 43496 47608 43502 47660
rect 64690 47648 64696 47660
rect 64651 47620 64696 47648
rect 64690 47608 64696 47620
rect 64748 47608 64754 47660
rect 4062 47540 4068 47592
rect 4120 47580 4126 47592
rect 43901 47583 43959 47589
rect 43901 47580 43913 47583
rect 4120 47552 43913 47580
rect 4120 47540 4126 47552
rect 43901 47549 43913 47552
rect 43947 47549 43959 47583
rect 65334 47580 65340 47592
rect 65295 47552 65340 47580
rect 43901 47543 43959 47549
rect 65334 47540 65340 47552
rect 65392 47540 65398 47592
rect 67174 47580 67180 47592
rect 67135 47552 67180 47580
rect 67174 47540 67180 47552
rect 67232 47540 67238 47592
rect 1104 47354 68816 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 68816 47354
rect 1104 47280 68816 47302
rect 65334 47200 65340 47252
rect 65392 47240 65398 47252
rect 65797 47243 65855 47249
rect 65797 47240 65809 47243
rect 65392 47212 65809 47240
rect 65392 47200 65398 47212
rect 65797 47209 65809 47212
rect 65843 47209 65855 47243
rect 65797 47203 65855 47209
rect 43530 47064 43536 47116
rect 43588 47104 43594 47116
rect 43625 47107 43683 47113
rect 43625 47104 43637 47107
rect 43588 47076 43637 47104
rect 43588 47064 43594 47076
rect 43625 47073 43637 47076
rect 43671 47104 43683 47107
rect 43806 47104 43812 47116
rect 43671 47076 43812 47104
rect 43671 47073 43683 47076
rect 43625 47067 43683 47073
rect 43806 47064 43812 47076
rect 43864 47064 43870 47116
rect 43901 47107 43959 47113
rect 43901 47073 43913 47107
rect 43947 47104 43959 47107
rect 44174 47104 44180 47116
rect 43947 47076 44180 47104
rect 43947 47073 43959 47076
rect 43901 47067 43959 47073
rect 44174 47064 44180 47076
rect 44232 47064 44238 47116
rect 45370 47104 45376 47116
rect 45331 47076 45376 47104
rect 45370 47064 45376 47076
rect 45428 47104 45434 47116
rect 45428 47076 45554 47104
rect 45428 47064 45434 47076
rect 44192 47036 44220 47064
rect 45097 47039 45155 47045
rect 45097 47036 45109 47039
rect 44192 47008 45109 47036
rect 45097 47005 45109 47008
rect 45143 47005 45155 47039
rect 45097 46999 45155 47005
rect 45526 46968 45554 47076
rect 62942 46968 62948 46980
rect 45526 46940 62948 46968
rect 62942 46928 62948 46940
rect 63000 46928 63006 46980
rect 1104 46810 68816 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 68816 46810
rect 1104 46736 68816 46758
rect 1104 46266 68816 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 68816 46266
rect 1104 46192 68816 46214
rect 37274 45908 37280 45960
rect 37332 45948 37338 45960
rect 37369 45951 37427 45957
rect 37369 45948 37381 45951
rect 37332 45920 37381 45948
rect 37332 45908 37338 45920
rect 37369 45917 37381 45920
rect 37415 45917 37427 45951
rect 37369 45911 37427 45917
rect 1104 45722 68816 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 68816 45722
rect 1104 45648 68816 45670
rect 37274 45472 37280 45484
rect 37235 45444 37280 45472
rect 37274 45432 37280 45444
rect 37332 45432 37338 45484
rect 48774 45432 48780 45484
rect 48832 45472 48838 45484
rect 49510 45472 49516 45484
rect 48832 45444 49516 45472
rect 48832 45432 48838 45444
rect 49510 45432 49516 45444
rect 49568 45432 49574 45484
rect 37458 45404 37464 45416
rect 37419 45376 37464 45404
rect 37458 45364 37464 45376
rect 37516 45364 37522 45416
rect 38470 45404 38476 45416
rect 38431 45376 38476 45404
rect 38470 45364 38476 45376
rect 38528 45364 38534 45416
rect 47578 45296 47584 45348
rect 47636 45336 47642 45348
rect 49789 45339 49847 45345
rect 49789 45336 49801 45339
rect 47636 45308 49801 45336
rect 47636 45296 47642 45308
rect 49789 45305 49801 45308
rect 49835 45336 49847 45339
rect 67450 45336 67456 45348
rect 49835 45308 67456 45336
rect 49835 45305 49847 45308
rect 49789 45299 49847 45305
rect 67450 45296 67456 45308
rect 67508 45296 67514 45348
rect 14734 45228 14740 45280
rect 14792 45268 14798 45280
rect 14921 45271 14979 45277
rect 14921 45268 14933 45271
rect 14792 45240 14933 45268
rect 14792 45228 14798 45240
rect 14921 45237 14933 45240
rect 14967 45237 14979 45271
rect 14921 45231 14979 45237
rect 66254 45228 66260 45280
rect 66312 45268 66318 45280
rect 67637 45271 67695 45277
rect 67637 45268 67649 45271
rect 66312 45240 67649 45268
rect 66312 45228 66318 45240
rect 67637 45237 67649 45240
rect 67683 45237 67695 45271
rect 67637 45231 67695 45237
rect 1104 45178 68816 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 68816 45178
rect 1104 45104 68816 45126
rect 36909 45067 36967 45073
rect 36909 45033 36921 45067
rect 36955 45064 36967 45067
rect 37458 45064 37464 45076
rect 36955 45036 37464 45064
rect 36955 45033 36967 45036
rect 36909 45027 36967 45033
rect 37458 45024 37464 45036
rect 37516 45024 37522 45076
rect 3418 44956 3424 45008
rect 3476 44996 3482 45008
rect 3476 44968 15240 44996
rect 3476 44956 3482 44968
rect 14734 44928 14740 44940
rect 14695 44900 14740 44928
rect 14734 44888 14740 44900
rect 14792 44888 14798 44940
rect 15212 44937 15240 44968
rect 15197 44931 15255 44937
rect 15197 44897 15209 44931
rect 15243 44897 15255 44931
rect 66254 44928 66260 44940
rect 66215 44900 66260 44928
rect 15197 44891 15255 44897
rect 66254 44888 66260 44900
rect 66312 44888 66318 44940
rect 68094 44928 68100 44940
rect 68055 44900 68100 44928
rect 68094 44888 68100 44900
rect 68152 44888 68158 44940
rect 22186 44820 22192 44872
rect 22244 44860 22250 44872
rect 28534 44860 28540 44872
rect 22244 44832 28540 44860
rect 22244 44820 22250 44832
rect 28534 44820 28540 44832
rect 28592 44860 28598 44872
rect 36817 44863 36875 44869
rect 36817 44860 36829 44863
rect 28592 44832 36829 44860
rect 28592 44820 28598 44832
rect 36817 44829 36829 44832
rect 36863 44829 36875 44863
rect 36817 44823 36875 44829
rect 14921 44795 14979 44801
rect 14921 44761 14933 44795
rect 14967 44792 14979 44795
rect 15102 44792 15108 44804
rect 14967 44764 15108 44792
rect 14967 44761 14979 44764
rect 14921 44755 14979 44761
rect 15102 44752 15108 44764
rect 15160 44752 15166 44804
rect 66438 44792 66444 44804
rect 66399 44764 66444 44792
rect 66438 44752 66444 44764
rect 66496 44752 66502 44804
rect 1104 44634 68816 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 68816 44634
rect 1104 44560 68816 44582
rect 15102 44520 15108 44532
rect 15063 44492 15108 44520
rect 15102 44480 15108 44492
rect 15160 44480 15166 44532
rect 66438 44480 66444 44532
rect 66496 44520 66502 44532
rect 67545 44523 67603 44529
rect 67545 44520 67557 44523
rect 66496 44492 67557 44520
rect 66496 44480 66502 44492
rect 67545 44489 67557 44492
rect 67591 44489 67603 44523
rect 67545 44483 67603 44489
rect 13722 44344 13728 44396
rect 13780 44384 13786 44396
rect 15013 44387 15071 44393
rect 15013 44384 15025 44387
rect 13780 44356 15025 44384
rect 13780 44344 13786 44356
rect 15013 44353 15025 44356
rect 15059 44353 15071 44387
rect 37734 44384 37740 44396
rect 37695 44356 37740 44384
rect 15013 44347 15071 44353
rect 37734 44344 37740 44356
rect 37792 44344 37798 44396
rect 43806 44344 43812 44396
rect 43864 44384 43870 44396
rect 44085 44387 44143 44393
rect 44085 44384 44097 44387
rect 43864 44356 44097 44384
rect 43864 44344 43870 44356
rect 44085 44353 44097 44356
rect 44131 44353 44143 44387
rect 67450 44384 67456 44396
rect 67411 44356 67456 44384
rect 44085 44347 44143 44353
rect 67450 44344 67456 44356
rect 67508 44344 67514 44396
rect 37918 44276 37924 44328
rect 37976 44316 37982 44328
rect 38013 44319 38071 44325
rect 38013 44316 38025 44319
rect 37976 44288 38025 44316
rect 37976 44276 37982 44288
rect 38013 44285 38025 44288
rect 38059 44316 38071 44319
rect 52086 44316 52092 44328
rect 38059 44288 52092 44316
rect 38059 44285 38071 44288
rect 38013 44279 38071 44285
rect 52086 44276 52092 44288
rect 52144 44276 52150 44328
rect 44082 44140 44088 44192
rect 44140 44180 44146 44192
rect 44177 44183 44235 44189
rect 44177 44180 44189 44183
rect 44140 44152 44189 44180
rect 44140 44140 44146 44152
rect 44177 44149 44189 44152
rect 44223 44180 44235 44183
rect 48774 44180 48780 44192
rect 44223 44152 48780 44180
rect 44223 44149 44235 44152
rect 44177 44143 44235 44149
rect 48774 44140 48780 44152
rect 48832 44140 48838 44192
rect 1104 44090 68816 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 68816 44090
rect 1104 44016 68816 44038
rect 52086 43772 52092 43784
rect 52047 43744 52092 43772
rect 52086 43732 52092 43744
rect 52144 43732 52150 43784
rect 52730 43772 52736 43784
rect 52691 43744 52736 43772
rect 52730 43732 52736 43744
rect 52788 43732 52794 43784
rect 52181 43707 52239 43713
rect 52181 43673 52193 43707
rect 52227 43704 52239 43707
rect 52917 43707 52975 43713
rect 52917 43704 52929 43707
rect 52227 43676 52929 43704
rect 52227 43673 52239 43676
rect 52181 43667 52239 43673
rect 52917 43673 52929 43676
rect 52963 43673 52975 43707
rect 52917 43667 52975 43673
rect 54573 43707 54631 43713
rect 54573 43673 54585 43707
rect 54619 43704 54631 43707
rect 66162 43704 66168 43716
rect 54619 43676 66168 43704
rect 54619 43673 54631 43676
rect 54573 43667 54631 43673
rect 66162 43664 66168 43676
rect 66220 43664 66226 43716
rect 1104 43546 68816 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 68816 43546
rect 1104 43472 68816 43494
rect 52730 43256 52736 43308
rect 52788 43296 52794 43308
rect 53009 43299 53067 43305
rect 53009 43296 53021 43299
rect 52788 43268 53021 43296
rect 52788 43256 52794 43268
rect 53009 43265 53021 43268
rect 53055 43265 53067 43299
rect 53009 43259 53067 43265
rect 1104 43002 68816 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 68816 43002
rect 1104 42928 68816 42950
rect 52086 42644 52092 42696
rect 52144 42684 52150 42696
rect 54481 42687 54539 42693
rect 54481 42684 54493 42687
rect 52144 42656 54493 42684
rect 52144 42644 52150 42656
rect 54481 42653 54493 42656
rect 54527 42653 54539 42687
rect 54481 42647 54539 42653
rect 54573 42551 54631 42557
rect 54573 42517 54585 42551
rect 54619 42548 54631 42551
rect 54938 42548 54944 42560
rect 54619 42520 54944 42548
rect 54619 42517 54631 42520
rect 54573 42511 54631 42517
rect 54938 42508 54944 42520
rect 54996 42508 55002 42560
rect 1104 42458 68816 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 68816 42458
rect 1104 42384 68816 42406
rect 54938 42276 54944 42288
rect 54899 42248 54944 42276
rect 54938 42236 54944 42248
rect 54996 42236 55002 42288
rect 12618 42168 12624 42220
rect 12676 42208 12682 42220
rect 13722 42208 13728 42220
rect 12676 42180 13728 42208
rect 12676 42168 12682 42180
rect 13722 42168 13728 42180
rect 13780 42208 13786 42220
rect 19981 42211 20039 42217
rect 19981 42208 19993 42211
rect 13780 42180 19993 42208
rect 13780 42168 13786 42180
rect 19981 42177 19993 42180
rect 20027 42208 20039 42211
rect 44082 42208 44088 42220
rect 20027 42180 26234 42208
rect 44043 42180 44088 42208
rect 20027 42177 20039 42180
rect 19981 42171 20039 42177
rect 20622 42100 20628 42152
rect 20680 42140 20686 42152
rect 20809 42143 20867 42149
rect 20809 42140 20821 42143
rect 20680 42112 20821 42140
rect 20680 42100 20686 42112
rect 20809 42109 20821 42112
rect 20855 42140 20867 42143
rect 24854 42140 24860 42152
rect 20855 42112 24860 42140
rect 20855 42109 20867 42112
rect 20809 42103 20867 42109
rect 24854 42100 24860 42112
rect 24912 42100 24918 42152
rect 26206 42140 26234 42180
rect 44082 42168 44088 42180
rect 44140 42168 44146 42220
rect 37734 42140 37740 42152
rect 26206 42112 37740 42140
rect 37734 42100 37740 42112
rect 37792 42140 37798 42152
rect 43530 42140 43536 42152
rect 37792 42112 43536 42140
rect 37792 42100 37798 42112
rect 43530 42100 43536 42112
rect 43588 42140 43594 42152
rect 44269 42143 44327 42149
rect 44269 42140 44281 42143
rect 43588 42112 44281 42140
rect 43588 42100 43594 42112
rect 44269 42109 44281 42112
rect 44315 42109 44327 42143
rect 44269 42103 44327 42109
rect 54297 42143 54355 42149
rect 54297 42109 54309 42143
rect 54343 42140 54355 42143
rect 54757 42143 54815 42149
rect 54757 42140 54769 42143
rect 54343 42112 54769 42140
rect 54343 42109 54355 42112
rect 54297 42103 54355 42109
rect 54757 42109 54769 42112
rect 54803 42109 54815 42143
rect 56502 42140 56508 42152
rect 56463 42112 56508 42140
rect 54757 42103 54815 42109
rect 56502 42100 56508 42112
rect 56560 42100 56566 42152
rect 1104 41914 68816 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 68816 41914
rect 1104 41840 68816 41862
rect 24854 41420 24860 41472
rect 24912 41460 24918 41472
rect 26418 41460 26424 41472
rect 24912 41432 26424 41460
rect 24912 41420 24918 41432
rect 26418 41420 26424 41432
rect 26476 41420 26482 41472
rect 1104 41370 68816 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 68816 41370
rect 1104 41296 68816 41318
rect 57241 41191 57299 41197
rect 57241 41157 57253 41191
rect 57287 41188 57299 41191
rect 58069 41191 58127 41197
rect 58069 41188 58081 41191
rect 57287 41160 58081 41188
rect 57287 41157 57299 41160
rect 57241 41151 57299 41157
rect 58069 41157 58081 41160
rect 58115 41157 58127 41191
rect 58069 41151 58127 41157
rect 44358 41080 44364 41132
rect 44416 41120 44422 41132
rect 57149 41123 57207 41129
rect 57149 41120 57161 41123
rect 44416 41092 57161 41120
rect 44416 41080 44422 41092
rect 57149 41089 57161 41092
rect 57195 41089 57207 41123
rect 57149 41083 57207 41089
rect 57882 41052 57888 41064
rect 57843 41024 57888 41052
rect 57882 41012 57888 41024
rect 57940 41012 57946 41064
rect 59725 41055 59783 41061
rect 59725 41021 59737 41055
rect 59771 41052 59783 41055
rect 66162 41052 66168 41064
rect 59771 41024 66168 41052
rect 59771 41021 59783 41024
rect 59725 41015 59783 41021
rect 66162 41012 66168 41024
rect 66220 41012 66226 41064
rect 1104 40826 68816 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 68816 40826
rect 1104 40752 68816 40774
rect 57882 40712 57888 40724
rect 57843 40684 57888 40712
rect 57882 40672 57888 40684
rect 57940 40672 57946 40724
rect 1104 40282 68816 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 68816 40282
rect 1104 40208 68816 40230
rect 3050 40060 3056 40112
rect 3108 40100 3114 40112
rect 23842 40100 23848 40112
rect 3108 40072 23848 40100
rect 3108 40060 3114 40072
rect 23842 40060 23848 40072
rect 23900 40060 23906 40112
rect 9582 39788 9588 39840
rect 9640 39828 9646 39840
rect 9769 39831 9827 39837
rect 9769 39828 9781 39831
rect 9640 39800 9781 39828
rect 9640 39788 9646 39800
rect 9769 39797 9781 39800
rect 9815 39797 9827 39831
rect 35342 39828 35348 39840
rect 35303 39800 35348 39828
rect 9769 39791 9827 39797
rect 35342 39788 35348 39800
rect 35400 39788 35406 39840
rect 60458 39788 60464 39840
rect 60516 39828 60522 39840
rect 60737 39831 60795 39837
rect 60737 39828 60749 39831
rect 60516 39800 60749 39828
rect 60516 39788 60522 39800
rect 60737 39797 60749 39800
rect 60783 39797 60795 39831
rect 60737 39791 60795 39797
rect 63218 39788 63224 39840
rect 63276 39828 63282 39840
rect 63865 39831 63923 39837
rect 63865 39828 63877 39831
rect 63276 39800 63877 39828
rect 63276 39788 63282 39800
rect 63865 39797 63877 39800
rect 63911 39797 63923 39831
rect 63865 39791 63923 39797
rect 1104 39738 68816 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 68816 39738
rect 1104 39664 68816 39686
rect 6886 39528 10088 39556
rect 3326 39312 3332 39364
rect 3384 39352 3390 39364
rect 6886 39352 6914 39528
rect 9582 39488 9588 39500
rect 9543 39460 9588 39488
rect 9582 39448 9588 39460
rect 9640 39448 9646 39500
rect 10060 39497 10088 39528
rect 10045 39491 10103 39497
rect 10045 39457 10057 39491
rect 10091 39457 10103 39491
rect 10045 39451 10103 39457
rect 22094 39448 22100 39500
rect 22152 39488 22158 39500
rect 23109 39491 23167 39497
rect 23109 39488 23121 39491
rect 22152 39460 23121 39488
rect 22152 39448 22158 39460
rect 23109 39457 23121 39460
rect 23155 39457 23167 39491
rect 23109 39451 23167 39457
rect 35069 39491 35127 39497
rect 35069 39457 35081 39491
rect 35115 39488 35127 39491
rect 35342 39488 35348 39500
rect 35115 39460 35348 39488
rect 35115 39457 35127 39460
rect 35069 39451 35127 39457
rect 35342 39448 35348 39460
rect 35400 39448 35406 39500
rect 36906 39488 36912 39500
rect 36867 39460 36912 39488
rect 36906 39448 36912 39460
rect 36964 39448 36970 39500
rect 60458 39488 60464 39500
rect 60419 39460 60464 39488
rect 60458 39448 60464 39460
rect 60516 39448 60522 39500
rect 62022 39488 62028 39500
rect 61983 39460 62028 39488
rect 62022 39448 62028 39460
rect 62080 39448 62086 39500
rect 63218 39488 63224 39500
rect 63179 39460 63224 39488
rect 63218 39448 63224 39460
rect 63276 39448 63282 39500
rect 64782 39488 64788 39500
rect 64743 39460 64788 39488
rect 64782 39448 64788 39460
rect 64840 39448 64846 39500
rect 22278 39380 22284 39432
rect 22336 39420 22342 39432
rect 22465 39423 22523 39429
rect 22465 39420 22477 39423
rect 22336 39392 22477 39420
rect 22336 39380 22342 39392
rect 22465 39389 22477 39392
rect 22511 39389 22523 39423
rect 22465 39383 22523 39389
rect 3384 39324 6914 39352
rect 9769 39355 9827 39361
rect 3384 39312 3390 39324
rect 9769 39321 9781 39355
rect 9815 39352 9827 39355
rect 9858 39352 9864 39364
rect 9815 39324 9864 39352
rect 9815 39321 9827 39324
rect 9769 39315 9827 39321
rect 9858 39312 9864 39324
rect 9916 39312 9922 39364
rect 34882 39312 34888 39364
rect 34940 39352 34946 39364
rect 35253 39355 35311 39361
rect 35253 39352 35265 39355
rect 34940 39324 35265 39352
rect 34940 39312 34946 39324
rect 35253 39321 35265 39324
rect 35299 39321 35311 39355
rect 60642 39352 60648 39364
rect 60603 39324 60648 39352
rect 35253 39315 35311 39321
rect 60642 39312 60648 39324
rect 60700 39312 60706 39364
rect 63405 39355 63463 39361
rect 63405 39321 63417 39355
rect 63451 39352 63463 39355
rect 63494 39352 63500 39364
rect 63451 39324 63500 39352
rect 63451 39321 63463 39324
rect 63405 39315 63463 39321
rect 63494 39312 63500 39324
rect 63552 39312 63558 39364
rect 1104 39194 68816 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 68816 39194
rect 1104 39120 68816 39142
rect 9858 39080 9864 39092
rect 9819 39052 9864 39080
rect 9858 39040 9864 39052
rect 9916 39040 9922 39092
rect 34882 39080 34888 39092
rect 34843 39052 34888 39080
rect 34882 39040 34888 39052
rect 34940 39040 34946 39092
rect 60461 39083 60519 39089
rect 60461 39049 60473 39083
rect 60507 39080 60519 39083
rect 60642 39080 60648 39092
rect 60507 39052 60648 39080
rect 60507 39049 60519 39052
rect 60461 39043 60519 39049
rect 60642 39040 60648 39052
rect 60700 39040 60706 39092
rect 63494 39080 63500 39092
rect 63455 39052 63500 39080
rect 63494 39040 63500 39052
rect 63552 39040 63558 39092
rect 24118 39012 24124 39024
rect 24079 38984 24124 39012
rect 24118 38972 24124 38984
rect 24176 38972 24182 39024
rect 48774 39012 48780 39024
rect 47688 38984 48780 39012
rect 9766 38944 9772 38956
rect 9727 38916 9772 38944
rect 9766 38904 9772 38916
rect 9824 38904 9830 38956
rect 22278 38944 22284 38956
rect 22239 38916 22284 38944
rect 22278 38904 22284 38916
rect 22336 38904 22342 38956
rect 34698 38904 34704 38956
rect 34756 38944 34762 38956
rect 34793 38947 34851 38953
rect 34793 38944 34805 38947
rect 34756 38916 34805 38944
rect 34756 38904 34762 38916
rect 34793 38913 34805 38916
rect 34839 38913 34851 38947
rect 34793 38907 34851 38913
rect 44358 38904 44364 38956
rect 44416 38944 44422 38956
rect 47688 38953 47716 38984
rect 48774 38972 48780 38984
rect 48832 38972 48838 39024
rect 44637 38947 44695 38953
rect 44637 38944 44649 38947
rect 44416 38916 44649 38944
rect 44416 38904 44422 38916
rect 44637 38913 44649 38916
rect 44683 38913 44695 38947
rect 44637 38907 44695 38913
rect 47673 38947 47731 38953
rect 47673 38913 47685 38947
rect 47719 38913 47731 38947
rect 47673 38907 47731 38913
rect 47949 38947 48007 38953
rect 47949 38913 47961 38947
rect 47995 38944 48007 38947
rect 60369 38947 60427 38953
rect 60369 38944 60381 38947
rect 47995 38916 60381 38944
rect 47995 38913 48007 38916
rect 47949 38907 48007 38913
rect 60369 38913 60381 38916
rect 60415 38944 60427 38947
rect 61838 38944 61844 38956
rect 60415 38916 61844 38944
rect 60415 38913 60427 38916
rect 60369 38907 60427 38913
rect 22462 38876 22468 38888
rect 22423 38848 22468 38876
rect 22462 38836 22468 38848
rect 22520 38836 22526 38888
rect 46382 38836 46388 38888
rect 46440 38876 46446 38888
rect 47964 38876 47992 38907
rect 61838 38904 61844 38916
rect 61896 38904 61902 38956
rect 63402 38944 63408 38956
rect 63363 38916 63408 38944
rect 63402 38904 63408 38916
rect 63460 38904 63466 38956
rect 46440 38848 47992 38876
rect 46440 38836 46446 38848
rect 44729 38743 44787 38749
rect 44729 38709 44741 38743
rect 44775 38740 44787 38743
rect 45186 38740 45192 38752
rect 44775 38712 45192 38740
rect 44775 38709 44787 38712
rect 44729 38703 44787 38709
rect 45186 38700 45192 38712
rect 45244 38700 45250 38752
rect 1104 38650 68816 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 68816 38650
rect 1104 38576 68816 38598
rect 21453 38539 21511 38545
rect 21453 38505 21465 38539
rect 21499 38536 21511 38539
rect 22462 38536 22468 38548
rect 21499 38508 22468 38536
rect 21499 38505 21511 38508
rect 21453 38499 21511 38505
rect 22462 38496 22468 38508
rect 22520 38496 22526 38548
rect 3418 38360 3424 38412
rect 3476 38400 3482 38412
rect 32769 38403 32827 38409
rect 32769 38400 32781 38403
rect 3476 38372 32781 38400
rect 3476 38360 3482 38372
rect 32769 38369 32781 38372
rect 32815 38369 32827 38403
rect 45186 38400 45192 38412
rect 45147 38372 45192 38400
rect 32769 38363 32827 38369
rect 45186 38360 45192 38372
rect 45244 38360 45250 38412
rect 21358 38332 21364 38344
rect 21319 38304 21364 38332
rect 21358 38292 21364 38304
rect 21416 38292 21422 38344
rect 22002 38332 22008 38344
rect 21963 38304 22008 38332
rect 22002 38292 22008 38304
rect 22060 38292 22066 38344
rect 23842 38332 23848 38344
rect 23803 38304 23848 38332
rect 23842 38292 23848 38304
rect 23900 38292 23906 38344
rect 32306 38332 32312 38344
rect 32267 38304 32312 38332
rect 32306 38292 32312 38304
rect 32364 38292 32370 38344
rect 44453 38335 44511 38341
rect 44453 38301 44465 38335
rect 44499 38332 44511 38335
rect 45005 38335 45063 38341
rect 45005 38332 45017 38335
rect 44499 38304 45017 38332
rect 44499 38301 44511 38304
rect 44453 38295 44511 38301
rect 45005 38301 45017 38304
rect 45051 38301 45063 38335
rect 51534 38332 51540 38344
rect 51495 38304 51540 38332
rect 45005 38295 45063 38301
rect 51534 38292 51540 38304
rect 51592 38292 51598 38344
rect 22189 38267 22247 38273
rect 22189 38233 22201 38267
rect 22235 38264 22247 38267
rect 22646 38264 22652 38276
rect 22235 38236 22652 38264
rect 22235 38233 22247 38236
rect 22189 38227 22247 38233
rect 22646 38224 22652 38236
rect 22704 38224 22710 38276
rect 32493 38267 32551 38273
rect 32493 38233 32505 38267
rect 32539 38264 32551 38267
rect 33502 38264 33508 38276
rect 32539 38236 33508 38264
rect 32539 38233 32551 38236
rect 32493 38227 32551 38233
rect 33502 38224 33508 38236
rect 33560 38224 33566 38276
rect 46842 38264 46848 38276
rect 46803 38236 46848 38264
rect 46842 38224 46848 38236
rect 46900 38224 46906 38276
rect 1104 38106 68816 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 68816 38106
rect 1104 38032 68816 38054
rect 22646 37992 22652 38004
rect 22607 37964 22652 37992
rect 22646 37952 22652 37964
rect 22704 37952 22710 38004
rect 33502 37992 33508 38004
rect 33463 37964 33508 37992
rect 33502 37952 33508 37964
rect 33560 37952 33566 38004
rect 7190 37924 7196 37936
rect 6886 37896 7196 37924
rect 6641 37859 6699 37865
rect 6641 37825 6653 37859
rect 6687 37856 6699 37859
rect 6886 37856 6914 37896
rect 7190 37884 7196 37896
rect 7248 37924 7254 37936
rect 20809 37927 20867 37933
rect 20809 37924 20821 37927
rect 7248 37896 20821 37924
rect 7248 37884 7254 37896
rect 20809 37893 20821 37896
rect 20855 37924 20867 37927
rect 28718 37924 28724 37936
rect 20855 37896 28724 37924
rect 20855 37893 20867 37896
rect 20809 37887 20867 37893
rect 28718 37884 28724 37896
rect 28776 37884 28782 37936
rect 6687 37828 6914 37856
rect 20533 37859 20591 37865
rect 6687 37825 6699 37828
rect 6641 37819 6699 37825
rect 20533 37825 20545 37859
rect 20579 37856 20591 37859
rect 20622 37856 20628 37868
rect 20579 37828 20628 37856
rect 20579 37825 20591 37828
rect 20533 37819 20591 37825
rect 20622 37816 20628 37828
rect 20680 37816 20686 37868
rect 22554 37856 22560 37868
rect 22515 37828 22560 37856
rect 22554 37816 22560 37828
rect 22612 37816 22618 37868
rect 32306 37816 32312 37868
rect 32364 37856 32370 37868
rect 32953 37859 33011 37865
rect 32953 37856 32965 37859
rect 32364 37828 32965 37856
rect 32364 37816 32370 37828
rect 32953 37825 32965 37828
rect 32999 37825 33011 37859
rect 32953 37819 33011 37825
rect 33413 37859 33471 37865
rect 33413 37825 33425 37859
rect 33459 37856 33471 37859
rect 46382 37856 46388 37868
rect 33459 37828 46388 37856
rect 33459 37825 33471 37828
rect 33413 37819 33471 37825
rect 28810 37748 28816 37800
rect 28868 37788 28874 37800
rect 33428 37788 33456 37819
rect 46382 37816 46388 37828
rect 46440 37816 46446 37868
rect 48774 37856 48780 37868
rect 48735 37828 48780 37856
rect 48774 37816 48780 37828
rect 48832 37816 48838 37868
rect 51166 37856 51172 37868
rect 51127 37828 51172 37856
rect 51166 37816 51172 37828
rect 51224 37816 51230 37868
rect 28868 37760 33456 37788
rect 28868 37748 28874 37760
rect 48958 37748 48964 37800
rect 49016 37788 49022 37800
rect 49053 37791 49111 37797
rect 49053 37788 49065 37791
rect 49016 37760 49065 37788
rect 49016 37748 49022 37760
rect 49053 37757 49065 37760
rect 49099 37788 49111 37791
rect 63402 37788 63408 37800
rect 49099 37760 63408 37788
rect 49099 37757 49111 37760
rect 49053 37751 49111 37757
rect 63402 37748 63408 37760
rect 63460 37748 63466 37800
rect 6546 37612 6552 37664
rect 6604 37652 6610 37664
rect 6733 37655 6791 37661
rect 6733 37652 6745 37655
rect 6604 37624 6745 37652
rect 6604 37612 6610 37624
rect 6733 37621 6745 37624
rect 6779 37621 6791 37655
rect 51258 37652 51264 37664
rect 51219 37624 51264 37652
rect 6733 37615 6791 37621
rect 51258 37612 51264 37624
rect 51316 37612 51322 37664
rect 1104 37562 68816 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 68816 37562
rect 1104 37488 68816 37510
rect 4982 37272 4988 37324
rect 5040 37312 5046 37324
rect 20073 37315 20131 37321
rect 20073 37312 20085 37315
rect 5040 37284 20085 37312
rect 5040 37272 5046 37284
rect 20073 37281 20085 37284
rect 20119 37312 20131 37315
rect 21358 37312 21364 37324
rect 20119 37284 21364 37312
rect 20119 37281 20131 37284
rect 20073 37275 20131 37281
rect 21358 37272 21364 37284
rect 21416 37272 21422 37324
rect 51353 37315 51411 37321
rect 51353 37281 51365 37315
rect 51399 37312 51411 37315
rect 51534 37312 51540 37324
rect 51399 37284 51540 37312
rect 51399 37281 51411 37284
rect 51353 37275 51411 37281
rect 51534 37272 51540 37284
rect 51592 37272 51598 37324
rect 5258 37204 5264 37256
rect 5316 37244 5322 37256
rect 5445 37247 5503 37253
rect 5445 37244 5457 37247
rect 5316 37216 5457 37244
rect 5316 37204 5322 37216
rect 5445 37213 5457 37216
rect 5491 37213 5503 37247
rect 5445 37207 5503 37213
rect 6362 37204 6368 37256
rect 6420 37244 6426 37256
rect 6457 37247 6515 37253
rect 6457 37244 6469 37247
rect 6420 37216 6469 37244
rect 6420 37204 6426 37216
rect 6457 37213 6469 37216
rect 6503 37213 6515 37247
rect 6457 37207 6515 37213
rect 19797 37247 19855 37253
rect 19797 37213 19809 37247
rect 19843 37244 19855 37247
rect 20622 37244 20628 37256
rect 19843 37216 20628 37244
rect 19843 37213 19855 37216
rect 19797 37207 19855 37213
rect 20622 37204 20628 37216
rect 20680 37244 20686 37256
rect 21545 37247 21603 37253
rect 21545 37244 21557 37247
rect 20680 37216 21557 37244
rect 20680 37204 20686 37216
rect 21545 37213 21557 37216
rect 21591 37213 21603 37247
rect 21545 37207 21603 37213
rect 21821 37247 21879 37253
rect 21821 37213 21833 37247
rect 21867 37244 21879 37247
rect 22186 37244 22192 37256
rect 21867 37216 22192 37244
rect 21867 37213 21879 37216
rect 21821 37207 21879 37213
rect 22186 37204 22192 37216
rect 22244 37204 22250 37256
rect 53193 37247 53251 37253
rect 53193 37213 53205 37247
rect 53239 37244 53251 37247
rect 53374 37244 53380 37256
rect 53239 37216 53380 37244
rect 53239 37213 53251 37216
rect 53193 37207 53251 37213
rect 53374 37204 53380 37216
rect 53432 37204 53438 37256
rect 20898 37176 20904 37188
rect 20859 37148 20904 37176
rect 20898 37136 20904 37148
rect 20956 37176 20962 37188
rect 35434 37176 35440 37188
rect 20956 37148 35440 37176
rect 20956 37136 20962 37148
rect 35434 37136 35440 37148
rect 35492 37136 35498 37188
rect 51258 37136 51264 37188
rect 51316 37176 51322 37188
rect 51537 37179 51595 37185
rect 51537 37176 51549 37179
rect 51316 37148 51549 37176
rect 51316 37136 51322 37148
rect 51537 37145 51549 37148
rect 51583 37145 51595 37179
rect 51537 37139 51595 37145
rect 1104 37018 68816 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 68816 37018
rect 1104 36944 68816 36966
rect 6546 36836 6552 36848
rect 6507 36808 6552 36836
rect 6546 36796 6552 36808
rect 6604 36796 6610 36848
rect 4982 36728 4988 36780
rect 5040 36768 5046 36780
rect 5445 36771 5503 36777
rect 5445 36768 5457 36771
rect 5040 36740 5457 36768
rect 5040 36728 5046 36740
rect 5445 36737 5457 36740
rect 5491 36737 5503 36771
rect 6362 36768 6368 36780
rect 6323 36740 6368 36768
rect 5445 36731 5503 36737
rect 6362 36728 6368 36740
rect 6420 36728 6426 36780
rect 20622 36768 20628 36780
rect 20583 36740 20628 36768
rect 20622 36728 20628 36740
rect 20680 36728 20686 36780
rect 38838 36768 38844 36780
rect 38751 36740 38844 36768
rect 38838 36728 38844 36740
rect 38896 36768 38902 36780
rect 43898 36768 43904 36780
rect 38896 36740 43904 36768
rect 38896 36728 38902 36740
rect 43898 36728 43904 36740
rect 43956 36728 43962 36780
rect 4614 36660 4620 36712
rect 4672 36700 4678 36712
rect 6825 36703 6883 36709
rect 6825 36700 6837 36703
rect 4672 36672 6837 36700
rect 4672 36660 4678 36672
rect 6825 36669 6837 36672
rect 6871 36669 6883 36703
rect 6825 36663 6883 36669
rect 9766 36660 9772 36712
rect 9824 36700 9830 36712
rect 20901 36703 20959 36709
rect 20901 36700 20913 36703
rect 9824 36672 20913 36700
rect 9824 36660 9830 36672
rect 20901 36669 20913 36672
rect 20947 36700 20959 36703
rect 34698 36700 34704 36712
rect 20947 36672 34704 36700
rect 20947 36669 20959 36672
rect 20901 36663 20959 36669
rect 34698 36660 34704 36672
rect 34756 36660 34762 36712
rect 5442 36524 5448 36576
rect 5500 36564 5506 36576
rect 5537 36567 5595 36573
rect 5537 36564 5549 36567
rect 5500 36536 5549 36564
rect 5500 36524 5506 36536
rect 5537 36533 5549 36536
rect 5583 36533 5595 36567
rect 5537 36527 5595 36533
rect 38102 36524 38108 36576
rect 38160 36564 38166 36576
rect 38381 36567 38439 36573
rect 38381 36564 38393 36567
rect 38160 36536 38393 36564
rect 38160 36524 38166 36536
rect 38381 36533 38393 36536
rect 38427 36533 38439 36567
rect 38930 36564 38936 36576
rect 38891 36536 38936 36564
rect 38381 36527 38439 36533
rect 38930 36524 38936 36536
rect 38988 36524 38994 36576
rect 1104 36474 68816 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 68816 36474
rect 1104 36400 68816 36422
rect 20533 36363 20591 36369
rect 20533 36329 20545 36363
rect 20579 36360 20591 36363
rect 20622 36360 20628 36372
rect 20579 36332 20628 36360
rect 20579 36329 20591 36332
rect 20533 36323 20591 36329
rect 20622 36320 20628 36332
rect 20680 36320 20686 36372
rect 2866 36252 2872 36304
rect 2924 36292 2930 36304
rect 2924 36264 5764 36292
rect 2924 36252 2930 36264
rect 5258 36224 5264 36236
rect 5219 36196 5264 36224
rect 5258 36184 5264 36196
rect 5316 36184 5322 36236
rect 5442 36224 5448 36236
rect 5403 36196 5448 36224
rect 5442 36184 5448 36196
rect 5500 36184 5506 36236
rect 5736 36233 5764 36264
rect 5721 36227 5779 36233
rect 5721 36193 5733 36227
rect 5767 36193 5779 36227
rect 5721 36187 5779 36193
rect 20717 36159 20775 36165
rect 20717 36125 20729 36159
rect 20763 36156 20775 36159
rect 31386 36156 31392 36168
rect 20763 36128 31392 36156
rect 20763 36125 20775 36128
rect 20717 36119 20775 36125
rect 31386 36116 31392 36128
rect 31444 36116 31450 36168
rect 1104 35930 68816 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 68816 35930
rect 1104 35856 68816 35878
rect 38838 35816 38844 35828
rect 37384 35788 38844 35816
rect 37384 35689 37412 35788
rect 38838 35776 38844 35788
rect 38896 35776 38902 35828
rect 38289 35751 38347 35757
rect 38289 35717 38301 35751
rect 38335 35748 38347 35751
rect 38930 35748 38936 35760
rect 38335 35720 38936 35748
rect 38335 35717 38347 35720
rect 38289 35711 38347 35717
rect 38930 35708 38936 35720
rect 38988 35708 38994 35760
rect 37369 35683 37427 35689
rect 37369 35649 37381 35683
rect 37415 35649 37427 35683
rect 38102 35680 38108 35692
rect 38063 35652 38108 35680
rect 37369 35643 37427 35649
rect 38102 35640 38108 35652
rect 38160 35640 38166 35692
rect 39758 35612 39764 35624
rect 39719 35584 39764 35612
rect 39758 35572 39764 35584
rect 39816 35572 39822 35624
rect 63034 35612 63040 35624
rect 62995 35584 63040 35612
rect 63034 35572 63040 35584
rect 63092 35572 63098 35624
rect 63221 35615 63279 35621
rect 63221 35581 63233 35615
rect 63267 35612 63279 35615
rect 63770 35612 63776 35624
rect 63267 35584 63776 35612
rect 63267 35581 63279 35584
rect 63221 35575 63279 35581
rect 63770 35572 63776 35584
rect 63828 35572 63834 35624
rect 64877 35615 64935 35621
rect 64877 35581 64889 35615
rect 64923 35612 64935 35615
rect 66070 35612 66076 35624
rect 64923 35584 66076 35612
rect 64923 35581 64935 35584
rect 64877 35575 64935 35581
rect 66070 35572 66076 35584
rect 66128 35572 66134 35624
rect 2774 35436 2780 35488
rect 2832 35476 2838 35488
rect 4614 35476 4620 35488
rect 2832 35448 4620 35476
rect 2832 35436 2838 35448
rect 4614 35436 4620 35448
rect 4672 35436 4678 35488
rect 37090 35436 37096 35488
rect 37148 35476 37154 35488
rect 37461 35479 37519 35485
rect 37461 35476 37473 35479
rect 37148 35448 37473 35476
rect 37148 35436 37154 35448
rect 37461 35445 37473 35448
rect 37507 35445 37519 35479
rect 37461 35439 37519 35445
rect 1104 35386 68816 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 68816 35386
rect 1104 35312 68816 35334
rect 63034 35232 63040 35284
rect 63092 35272 63098 35284
rect 63221 35275 63279 35281
rect 63221 35272 63233 35275
rect 63092 35244 63233 35272
rect 63092 35232 63098 35244
rect 63221 35241 63233 35244
rect 63267 35241 63279 35275
rect 63770 35272 63776 35284
rect 63731 35244 63776 35272
rect 63221 35235 63279 35241
rect 63770 35232 63776 35244
rect 63828 35232 63834 35284
rect 26206 35176 37412 35204
rect 3418 34892 3424 34944
rect 3476 34932 3482 34944
rect 26206 34932 26234 35176
rect 37090 35136 37096 35148
rect 37051 35108 37096 35136
rect 37090 35096 37096 35108
rect 37148 35096 37154 35148
rect 37384 35145 37412 35176
rect 37369 35139 37427 35145
rect 37369 35105 37381 35139
rect 37415 35105 37427 35139
rect 37369 35099 37427 35105
rect 36449 35071 36507 35077
rect 36449 35037 36461 35071
rect 36495 35068 36507 35071
rect 36909 35071 36967 35077
rect 36909 35068 36921 35071
rect 36495 35040 36921 35068
rect 36495 35037 36507 35040
rect 36449 35031 36507 35037
rect 36909 35037 36921 35040
rect 36955 35037 36967 35071
rect 63678 35068 63684 35080
rect 63639 35040 63684 35068
rect 36909 35031 36967 35037
rect 63678 35028 63684 35040
rect 63736 35028 63742 35080
rect 3476 34904 26234 34932
rect 3476 34892 3482 34904
rect 1104 34842 68816 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 68816 34842
rect 1104 34768 68816 34790
rect 1104 34298 68816 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 68816 34298
rect 1104 34224 68816 34246
rect 42334 33940 42340 33992
rect 42392 33980 42398 33992
rect 42429 33983 42487 33989
rect 42429 33980 42441 33983
rect 42392 33952 42441 33980
rect 42392 33940 42398 33952
rect 42429 33949 42441 33952
rect 42475 33949 42487 33983
rect 42429 33943 42487 33949
rect 42886 33940 42892 33992
rect 42944 33980 42950 33992
rect 43533 33983 43591 33989
rect 43533 33980 43545 33983
rect 42944 33952 43545 33980
rect 42944 33940 42950 33952
rect 43533 33949 43545 33952
rect 43579 33949 43591 33983
rect 43533 33943 43591 33949
rect 42702 33912 42708 33924
rect 42615 33884 42708 33912
rect 42702 33872 42708 33884
rect 42760 33912 42766 33924
rect 49050 33912 49056 33924
rect 42760 33884 49056 33912
rect 42760 33872 42766 33884
rect 49050 33872 49056 33884
rect 49108 33872 49114 33924
rect 1104 33754 68816 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 68816 33754
rect 1104 33680 68816 33702
rect 41417 33507 41475 33513
rect 41417 33473 41429 33507
rect 41463 33504 41475 33507
rect 42334 33504 42340 33516
rect 41463 33476 42340 33504
rect 41463 33473 41475 33476
rect 41417 33467 41475 33473
rect 42334 33464 42340 33476
rect 42392 33464 42398 33516
rect 42886 33504 42892 33516
rect 42847 33476 42892 33504
rect 42886 33464 42892 33476
rect 42944 33464 42950 33516
rect 67450 33504 67456 33516
rect 67411 33476 67456 33504
rect 67450 33464 67456 33476
rect 67508 33464 67514 33516
rect 41598 33436 41604 33448
rect 41559 33408 41604 33436
rect 41598 33396 41604 33408
rect 41656 33396 41662 33448
rect 43070 33436 43076 33448
rect 43031 33408 43076 33436
rect 43070 33396 43076 33408
rect 43128 33396 43134 33448
rect 44729 33439 44787 33445
rect 44729 33405 44741 33439
rect 44775 33436 44787 33439
rect 65518 33436 65524 33448
rect 44775 33408 65524 33436
rect 44775 33405 44787 33408
rect 44729 33399 44787 33405
rect 65518 33396 65524 33408
rect 65576 33396 65582 33448
rect 41616 33368 41644 33396
rect 44082 33368 44088 33380
rect 41616 33340 44088 33368
rect 44082 33328 44088 33340
rect 44140 33328 44146 33380
rect 62390 33300 62396 33312
rect 62351 33272 62396 33300
rect 62390 33260 62396 33272
rect 62448 33260 62454 33312
rect 66438 33260 66444 33312
rect 66496 33300 66502 33312
rect 67545 33303 67603 33309
rect 67545 33300 67557 33303
rect 66496 33272 67557 33300
rect 66496 33260 66502 33272
rect 67545 33269 67557 33272
rect 67591 33269 67603 33303
rect 67545 33263 67603 33269
rect 1104 33210 68816 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 68816 33210
rect 1104 33136 68816 33158
rect 43070 33056 43076 33108
rect 43128 33096 43134 33108
rect 43533 33099 43591 33105
rect 43533 33096 43545 33099
rect 43128 33068 43545 33096
rect 43128 33056 43134 33068
rect 43533 33065 43545 33068
rect 43579 33065 43591 33099
rect 51074 33096 51080 33108
rect 43533 33059 43591 33065
rect 45526 33068 51080 33096
rect 42153 32963 42211 32969
rect 42153 32929 42165 32963
rect 42199 32960 42211 32963
rect 43806 32960 43812 32972
rect 42199 32932 43812 32960
rect 42199 32929 42211 32932
rect 42153 32923 42211 32929
rect 43806 32920 43812 32932
rect 43864 32920 43870 32972
rect 42334 32852 42340 32904
rect 42392 32892 42398 32904
rect 42429 32895 42487 32901
rect 42429 32892 42441 32895
rect 42392 32864 42441 32892
rect 42392 32852 42398 32864
rect 42429 32861 42441 32864
rect 42475 32861 42487 32895
rect 42429 32855 42487 32861
rect 42978 32852 42984 32904
rect 43036 32892 43042 32904
rect 43441 32895 43499 32901
rect 43441 32892 43453 32895
rect 43036 32864 43453 32892
rect 43036 32852 43042 32864
rect 43441 32861 43453 32864
rect 43487 32861 43499 32895
rect 44082 32892 44088 32904
rect 44043 32864 44088 32892
rect 43441 32855 43499 32861
rect 44082 32852 44088 32864
rect 44140 32892 44146 32904
rect 45526 32892 45554 33068
rect 51074 33056 51080 33068
rect 51132 33096 51138 33108
rect 54202 33096 54208 33108
rect 51132 33068 54208 33096
rect 51132 33056 51138 33068
rect 54202 33056 54208 33068
rect 54260 33056 54266 33108
rect 62209 32963 62267 32969
rect 62209 32929 62221 32963
rect 62255 32960 62267 32963
rect 62390 32960 62396 32972
rect 62255 32932 62396 32960
rect 62255 32929 62267 32932
rect 62209 32923 62267 32929
rect 62390 32920 62396 32932
rect 62448 32920 62454 32972
rect 65794 32920 65800 32972
rect 65852 32960 65858 32972
rect 67913 32963 67971 32969
rect 67913 32960 67925 32963
rect 65852 32932 67925 32960
rect 65852 32920 65858 32932
rect 67913 32929 67925 32932
rect 67959 32929 67971 32963
rect 67913 32923 67971 32929
rect 44140 32864 45554 32892
rect 67085 32895 67143 32901
rect 44140 32852 44146 32864
rect 67085 32861 67097 32895
rect 67131 32892 67143 32895
rect 67450 32892 67456 32904
rect 67131 32864 67456 32892
rect 67131 32861 67143 32864
rect 67085 32855 67143 32861
rect 67450 32852 67456 32864
rect 67508 32852 67514 32904
rect 61930 32784 61936 32836
rect 61988 32824 61994 32836
rect 62393 32827 62451 32833
rect 62393 32824 62405 32827
rect 61988 32796 62405 32824
rect 61988 32784 61994 32796
rect 62393 32793 62405 32796
rect 62439 32793 62451 32827
rect 62393 32787 62451 32793
rect 64049 32827 64107 32833
rect 64049 32793 64061 32827
rect 64095 32824 64107 32827
rect 66162 32824 66168 32836
rect 64095 32796 66168 32824
rect 64095 32793 64107 32796
rect 64049 32787 64107 32793
rect 66162 32784 66168 32796
rect 66220 32784 66226 32836
rect 44082 32716 44088 32768
rect 44140 32756 44146 32768
rect 44177 32759 44235 32765
rect 44177 32756 44189 32759
rect 44140 32728 44189 32756
rect 44140 32716 44146 32728
rect 44177 32725 44189 32728
rect 44223 32725 44235 32759
rect 44177 32719 44235 32725
rect 65978 32716 65984 32768
rect 66036 32756 66042 32768
rect 67177 32759 67235 32765
rect 67177 32756 67189 32759
rect 66036 32728 67189 32756
rect 66036 32716 66042 32728
rect 67177 32725 67189 32728
rect 67223 32725 67235 32759
rect 67177 32719 67235 32725
rect 1104 32666 68816 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 68816 32666
rect 1104 32592 68816 32614
rect 61930 32552 61936 32564
rect 61891 32524 61936 32552
rect 61930 32512 61936 32524
rect 61988 32512 61994 32564
rect 37366 32444 37372 32496
rect 37424 32484 37430 32496
rect 42705 32487 42763 32493
rect 42705 32484 42717 32487
rect 37424 32456 42717 32484
rect 37424 32444 37430 32456
rect 42705 32453 42717 32456
rect 42751 32453 42763 32487
rect 44082 32484 44088 32496
rect 44043 32456 44088 32484
rect 42705 32447 42763 32453
rect 42334 32376 42340 32428
rect 42392 32416 42398 32428
rect 42429 32419 42487 32425
rect 42429 32416 42441 32419
rect 42392 32388 42441 32416
rect 42392 32376 42398 32388
rect 42429 32385 42441 32388
rect 42475 32385 42487 32419
rect 42429 32379 42487 32385
rect 42720 32280 42748 32447
rect 44082 32444 44088 32456
rect 44140 32444 44146 32496
rect 65978 32484 65984 32496
rect 65939 32456 65984 32484
rect 65978 32444 65984 32456
rect 66036 32444 66042 32496
rect 43806 32376 43812 32428
rect 43864 32416 43870 32428
rect 43901 32419 43959 32425
rect 43901 32416 43913 32419
rect 43864 32388 43913 32416
rect 43864 32376 43870 32388
rect 43901 32385 43913 32388
rect 43947 32385 43959 32419
rect 43901 32379 43959 32385
rect 60734 32376 60740 32428
rect 60792 32416 60798 32428
rect 61838 32416 61844 32428
rect 60792 32388 61844 32416
rect 60792 32376 60798 32388
rect 61838 32376 61844 32388
rect 61896 32376 61902 32428
rect 65794 32416 65800 32428
rect 65755 32388 65800 32416
rect 65794 32376 65800 32388
rect 65852 32376 65858 32428
rect 45462 32348 45468 32360
rect 45423 32320 45468 32348
rect 45462 32308 45468 32320
rect 45520 32308 45526 32360
rect 67542 32348 67548 32360
rect 67503 32320 67548 32348
rect 67542 32308 67548 32320
rect 67600 32308 67606 32360
rect 47578 32280 47584 32292
rect 42720 32252 47584 32280
rect 47578 32240 47584 32252
rect 47636 32240 47642 32292
rect 1104 32122 68816 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 68816 32122
rect 1104 32048 68816 32070
rect 66257 31875 66315 31881
rect 66257 31841 66269 31875
rect 66303 31872 66315 31875
rect 67634 31872 67640 31884
rect 66303 31844 67640 31872
rect 66303 31841 66315 31844
rect 66257 31835 66315 31841
rect 67634 31832 67640 31844
rect 67692 31832 67698 31884
rect 67818 31872 67824 31884
rect 67779 31844 67824 31872
rect 67818 31832 67824 31844
rect 67876 31832 67882 31884
rect 42337 31807 42395 31813
rect 42337 31773 42349 31807
rect 42383 31804 42395 31807
rect 42702 31804 42708 31816
rect 42383 31776 42708 31804
rect 42383 31773 42395 31776
rect 42337 31767 42395 31773
rect 42702 31764 42708 31776
rect 42760 31764 42766 31816
rect 66438 31736 66444 31748
rect 66399 31708 66444 31736
rect 66438 31696 66444 31708
rect 66496 31696 66502 31748
rect 42429 31671 42487 31677
rect 42429 31637 42441 31671
rect 42475 31668 42487 31671
rect 42610 31668 42616 31680
rect 42475 31640 42616 31668
rect 42475 31637 42487 31640
rect 42429 31631 42487 31637
rect 42610 31628 42616 31640
rect 42668 31628 42674 31680
rect 1104 31578 68816 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 68816 31578
rect 1104 31504 68816 31526
rect 42610 31396 42616 31408
rect 42571 31368 42616 31396
rect 42610 31356 42616 31368
rect 42668 31356 42674 31408
rect 59081 31399 59139 31405
rect 59081 31365 59093 31399
rect 59127 31396 59139 31399
rect 59817 31399 59875 31405
rect 59817 31396 59829 31399
rect 59127 31368 59829 31396
rect 59127 31365 59139 31368
rect 59081 31359 59139 31365
rect 59817 31365 59829 31368
rect 59863 31365 59875 31399
rect 59817 31359 59875 31365
rect 49050 31288 49056 31340
rect 49108 31328 49114 31340
rect 58989 31331 59047 31337
rect 58989 31328 59001 31331
rect 49108 31300 59001 31328
rect 49108 31288 49114 31300
rect 58989 31297 59001 31300
rect 59035 31297 59047 31331
rect 67634 31328 67640 31340
rect 67595 31300 67640 31328
rect 58989 31291 59047 31297
rect 67634 31288 67640 31300
rect 67692 31288 67698 31340
rect 198 31220 204 31272
rect 256 31260 262 31272
rect 41877 31263 41935 31269
rect 256 31232 26234 31260
rect 256 31220 262 31232
rect 26206 31192 26234 31232
rect 41877 31229 41889 31263
rect 41923 31260 41935 31263
rect 42429 31263 42487 31269
rect 42429 31260 42441 31263
rect 41923 31232 42441 31260
rect 41923 31229 41935 31232
rect 41877 31223 41935 31229
rect 42429 31229 42441 31232
rect 42475 31229 42487 31263
rect 42429 31223 42487 31229
rect 42889 31263 42947 31269
rect 42889 31229 42901 31263
rect 42935 31229 42947 31263
rect 42889 31223 42947 31229
rect 59633 31263 59691 31269
rect 59633 31229 59645 31263
rect 59679 31260 59691 31263
rect 59814 31260 59820 31272
rect 59679 31232 59820 31260
rect 59679 31229 59691 31232
rect 59633 31223 59691 31229
rect 42904 31192 42932 31223
rect 59814 31220 59820 31232
rect 59872 31220 59878 31272
rect 61473 31263 61531 31269
rect 61473 31229 61485 31263
rect 61519 31260 61531 31263
rect 63126 31260 63132 31272
rect 61519 31232 63132 31260
rect 61519 31229 61531 31232
rect 61473 31223 61531 31229
rect 63126 31220 63132 31232
rect 63184 31220 63190 31272
rect 26206 31164 42932 31192
rect 42794 31084 42800 31136
rect 42852 31124 42858 31136
rect 43346 31124 43352 31136
rect 42852 31096 43352 31124
rect 42852 31084 42858 31096
rect 43346 31084 43352 31096
rect 43404 31124 43410 31136
rect 51166 31124 51172 31136
rect 43404 31096 51172 31124
rect 43404 31084 43410 31096
rect 51166 31084 51172 31096
rect 51224 31084 51230 31136
rect 1104 31034 68816 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 68816 31034
rect 1104 30960 68816 30982
rect 59814 30920 59820 30932
rect 59775 30892 59820 30920
rect 59814 30880 59820 30892
rect 59872 30880 59878 30932
rect 22554 30744 22560 30796
rect 22612 30784 22618 30796
rect 22612 30756 35894 30784
rect 22612 30744 22618 30756
rect 20622 30676 20628 30728
rect 20680 30716 20686 30728
rect 26418 30716 26424 30728
rect 20680 30688 26424 30716
rect 20680 30676 20686 30688
rect 26418 30676 26424 30688
rect 26476 30676 26482 30728
rect 27062 30716 27068 30728
rect 27023 30688 27068 30716
rect 27062 30676 27068 30688
rect 27120 30676 27126 30728
rect 26513 30651 26571 30657
rect 26513 30617 26525 30651
rect 26559 30648 26571 30651
rect 27249 30651 27307 30657
rect 27249 30648 27261 30651
rect 26559 30620 27261 30648
rect 26559 30617 26571 30620
rect 26513 30611 26571 30617
rect 27249 30617 27261 30620
rect 27295 30617 27307 30651
rect 28902 30648 28908 30660
rect 28863 30620 28908 30648
rect 27249 30611 27307 30617
rect 28902 30608 28908 30620
rect 28960 30608 28966 30660
rect 35866 30648 35894 30756
rect 42334 30716 42340 30728
rect 42295 30688 42340 30716
rect 42334 30676 42340 30688
rect 42392 30676 42398 30728
rect 42613 30651 42671 30657
rect 42613 30648 42625 30651
rect 35866 30620 42625 30648
rect 42613 30617 42625 30620
rect 42659 30648 42671 30651
rect 42794 30648 42800 30660
rect 42659 30620 42800 30648
rect 42659 30617 42671 30620
rect 42613 30611 42671 30617
rect 42794 30608 42800 30620
rect 42852 30608 42858 30660
rect 1104 30490 68816 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 68816 30490
rect 1104 30416 68816 30438
rect 42334 30268 42340 30320
rect 42392 30308 42398 30320
rect 42889 30311 42947 30317
rect 42889 30308 42901 30311
rect 42392 30280 42901 30308
rect 42392 30268 42398 30280
rect 42889 30277 42901 30280
rect 42935 30277 42947 30311
rect 42889 30271 42947 30277
rect 27062 30200 27068 30252
rect 27120 30240 27126 30252
rect 27249 30243 27307 30249
rect 27249 30240 27261 30243
rect 27120 30212 27261 30240
rect 27120 30200 27126 30212
rect 27249 30209 27261 30212
rect 27295 30209 27307 30243
rect 27249 30203 27307 30209
rect 8018 30172 8024 30184
rect 7979 30144 8024 30172
rect 8018 30132 8024 30144
rect 8076 30132 8082 30184
rect 8205 30175 8263 30181
rect 8205 30141 8217 30175
rect 8251 30172 8263 30175
rect 9030 30172 9036 30184
rect 8251 30144 9036 30172
rect 8251 30141 8263 30144
rect 8205 30135 8263 30141
rect 9030 30132 9036 30144
rect 9088 30132 9094 30184
rect 9125 30175 9183 30181
rect 9125 30141 9137 30175
rect 9171 30141 9183 30175
rect 9125 30135 9183 30141
rect 4062 30064 4068 30116
rect 4120 30104 4126 30116
rect 9140 30104 9168 30135
rect 63126 30132 63132 30184
rect 63184 30172 63190 30184
rect 66162 30172 66168 30184
rect 63184 30144 66168 30172
rect 63184 30132 63190 30144
rect 66162 30132 66168 30144
rect 66220 30132 66226 30184
rect 4120 30076 9168 30104
rect 4120 30064 4126 30076
rect 42978 30036 42984 30048
rect 42939 30008 42984 30036
rect 42978 29996 42984 30008
rect 43036 29996 43042 30048
rect 1104 29946 68816 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 68816 29946
rect 1104 29872 68816 29894
rect 8018 29792 8024 29844
rect 8076 29832 8082 29844
rect 8205 29835 8263 29841
rect 8205 29832 8217 29835
rect 8076 29804 8217 29832
rect 8076 29792 8082 29804
rect 8205 29801 8217 29804
rect 8251 29801 8263 29835
rect 9030 29832 9036 29844
rect 8991 29804 9036 29832
rect 8205 29795 8263 29801
rect 9030 29792 9036 29804
rect 9088 29792 9094 29844
rect 3418 29656 3424 29708
rect 3476 29696 3482 29708
rect 6089 29699 6147 29705
rect 6089 29696 6101 29699
rect 3476 29668 6101 29696
rect 3476 29656 3482 29668
rect 6089 29665 6101 29668
rect 6135 29665 6147 29699
rect 20898 29696 20904 29708
rect 6089 29659 6147 29665
rect 16546 29668 20904 29696
rect 4985 29631 5043 29637
rect 4985 29597 4997 29631
rect 5031 29597 5043 29631
rect 5626 29628 5632 29640
rect 5587 29600 5632 29628
rect 4985 29591 5043 29597
rect 5000 29492 5028 29591
rect 5626 29588 5632 29600
rect 5684 29588 5690 29640
rect 8941 29631 8999 29637
rect 8941 29597 8953 29631
rect 8987 29628 8999 29631
rect 9766 29628 9772 29640
rect 8987 29600 9772 29628
rect 8987 29597 8999 29600
rect 8941 29591 8999 29597
rect 9766 29588 9772 29600
rect 9824 29628 9830 29640
rect 10778 29628 10784 29640
rect 9824 29600 10784 29628
rect 9824 29588 9830 29600
rect 10778 29588 10784 29600
rect 10836 29588 10842 29640
rect 12158 29588 12164 29640
rect 12216 29628 12222 29640
rect 12437 29631 12495 29637
rect 12437 29628 12449 29631
rect 12216 29600 12449 29628
rect 12216 29588 12222 29600
rect 12437 29597 12449 29600
rect 12483 29597 12495 29631
rect 12437 29591 12495 29597
rect 5077 29563 5135 29569
rect 5077 29529 5089 29563
rect 5123 29560 5135 29563
rect 5813 29563 5871 29569
rect 5813 29560 5825 29563
rect 5123 29532 5825 29560
rect 5123 29529 5135 29532
rect 5077 29523 5135 29529
rect 5813 29529 5825 29532
rect 5859 29529 5871 29563
rect 5813 29523 5871 29529
rect 5442 29492 5448 29504
rect 5000 29464 5448 29492
rect 5442 29452 5448 29464
rect 5500 29492 5506 29504
rect 16546 29492 16574 29668
rect 20898 29656 20904 29668
rect 20956 29656 20962 29708
rect 43622 29588 43628 29640
rect 43680 29628 43686 29640
rect 43901 29631 43959 29637
rect 43901 29628 43913 29631
rect 43680 29600 43913 29628
rect 43680 29588 43686 29600
rect 43901 29597 43913 29600
rect 43947 29597 43959 29631
rect 43901 29591 43959 29597
rect 5500 29464 16574 29492
rect 5500 29452 5506 29464
rect 1104 29402 68816 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 68816 29402
rect 1104 29328 68816 29350
rect 5626 29112 5632 29164
rect 5684 29152 5690 29164
rect 6549 29155 6607 29161
rect 6549 29152 6561 29155
rect 5684 29124 6561 29152
rect 5684 29112 5690 29124
rect 6549 29121 6561 29124
rect 6595 29121 6607 29155
rect 12158 29152 12164 29164
rect 12119 29124 12164 29152
rect 6549 29115 6607 29121
rect 12158 29112 12164 29124
rect 12216 29112 12222 29164
rect 43622 29152 43628 29164
rect 43583 29124 43628 29152
rect 43622 29112 43628 29124
rect 43680 29112 43686 29164
rect 12345 29087 12403 29093
rect 12345 29053 12357 29087
rect 12391 29084 12403 29087
rect 12710 29084 12716 29096
rect 12391 29056 12716 29084
rect 12391 29053 12403 29056
rect 12345 29047 12403 29053
rect 12710 29044 12716 29056
rect 12768 29044 12774 29096
rect 12802 29044 12808 29096
rect 12860 29084 12866 29096
rect 43806 29084 43812 29096
rect 12860 29056 12905 29084
rect 43767 29056 43812 29084
rect 12860 29044 12866 29056
rect 43806 29044 43812 29056
rect 43864 29044 43870 29096
rect 45186 29084 45192 29096
rect 45147 29056 45192 29084
rect 45186 29044 45192 29056
rect 45244 29044 45250 29096
rect 1104 28858 68816 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 68816 28858
rect 1104 28784 68816 28806
rect 12710 28744 12716 28756
rect 12671 28716 12716 28744
rect 12710 28704 12716 28716
rect 12768 28704 12774 28756
rect 43625 28747 43683 28753
rect 43625 28713 43637 28747
rect 43671 28744 43683 28747
rect 43806 28744 43812 28756
rect 43671 28716 43812 28744
rect 43671 28713 43683 28716
rect 43625 28707 43683 28713
rect 43806 28704 43812 28716
rect 43864 28704 43870 28756
rect 4982 28540 4988 28552
rect 4943 28512 4988 28540
rect 4982 28500 4988 28512
rect 5040 28500 5046 28552
rect 5442 28540 5448 28552
rect 5403 28512 5448 28540
rect 5442 28500 5448 28512
rect 5500 28500 5506 28552
rect 12618 28540 12624 28552
rect 12579 28512 12624 28540
rect 12618 28500 12624 28512
rect 12676 28500 12682 28552
rect 43530 28540 43536 28552
rect 43491 28512 43536 28540
rect 43530 28500 43536 28512
rect 43588 28500 43594 28552
rect 54202 28540 54208 28552
rect 54163 28512 54208 28540
rect 54202 28500 54208 28512
rect 54260 28500 54266 28552
rect 54754 28500 54760 28552
rect 54812 28540 54818 28552
rect 55309 28543 55367 28549
rect 55309 28540 55321 28543
rect 54812 28512 55321 28540
rect 54812 28500 54818 28512
rect 55309 28509 55321 28512
rect 55355 28509 55367 28543
rect 55309 28503 55367 28509
rect 54297 28475 54355 28481
rect 54297 28441 54309 28475
rect 54343 28472 54355 28475
rect 55493 28475 55551 28481
rect 55493 28472 55505 28475
rect 54343 28444 55505 28472
rect 54343 28441 54355 28444
rect 54297 28435 54355 28441
rect 55493 28441 55505 28444
rect 55539 28441 55551 28475
rect 55493 28435 55551 28441
rect 57149 28475 57207 28481
rect 57149 28441 57161 28475
rect 57195 28472 57207 28475
rect 65518 28472 65524 28484
rect 57195 28444 65524 28472
rect 57195 28441 57207 28444
rect 57149 28435 57207 28441
rect 65518 28432 65524 28444
rect 65576 28432 65582 28484
rect 5534 28404 5540 28416
rect 5495 28376 5540 28404
rect 5534 28364 5540 28376
rect 5592 28364 5598 28416
rect 1104 28314 68816 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 68816 28314
rect 1104 28240 68816 28262
rect 9493 28067 9551 28073
rect 9493 28033 9505 28067
rect 9539 28064 9551 28067
rect 20622 28064 20628 28076
rect 9539 28036 20628 28064
rect 9539 28033 9551 28036
rect 9493 28027 9551 28033
rect 20622 28024 20628 28036
rect 20680 28024 20686 28076
rect 26973 28067 27031 28073
rect 26973 28033 26985 28067
rect 27019 28064 27031 28067
rect 41598 28064 41604 28076
rect 27019 28036 41604 28064
rect 27019 28033 27031 28036
rect 26973 28027 27031 28033
rect 41598 28024 41604 28036
rect 41656 28024 41662 28076
rect 54754 28064 54760 28076
rect 54715 28036 54760 28064
rect 54754 28024 54760 28036
rect 54812 28024 54818 28076
rect 9398 27820 9404 27872
rect 9456 27860 9462 27872
rect 9585 27863 9643 27869
rect 9585 27860 9597 27863
rect 9456 27832 9597 27860
rect 9456 27820 9462 27832
rect 9585 27829 9597 27832
rect 9631 27829 9643 27863
rect 10318 27860 10324 27872
rect 10279 27832 10324 27860
rect 9585 27823 9643 27829
rect 10318 27820 10324 27832
rect 10376 27820 10382 27872
rect 26234 27820 26240 27872
rect 26292 27860 26298 27872
rect 27062 27860 27068 27872
rect 26292 27832 26337 27860
rect 27023 27832 27068 27860
rect 26292 27820 26298 27832
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 1104 27770 68816 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 68816 27770
rect 1104 27696 68816 27718
rect 3970 27548 3976 27600
rect 4028 27588 4034 27600
rect 10318 27588 10324 27600
rect 4028 27560 5672 27588
rect 4028 27548 4034 27560
rect 4982 27480 4988 27532
rect 5040 27520 5046 27532
rect 5077 27523 5135 27529
rect 5077 27520 5089 27523
rect 5040 27492 5089 27520
rect 5040 27480 5046 27492
rect 5077 27489 5089 27492
rect 5123 27489 5135 27523
rect 5077 27483 5135 27489
rect 5261 27523 5319 27529
rect 5261 27489 5273 27523
rect 5307 27520 5319 27523
rect 5534 27520 5540 27532
rect 5307 27492 5540 27520
rect 5307 27489 5319 27492
rect 5261 27483 5319 27489
rect 5534 27480 5540 27492
rect 5592 27480 5598 27532
rect 5644 27529 5672 27560
rect 9232 27560 10324 27588
rect 9232 27529 9260 27560
rect 10318 27548 10324 27560
rect 10376 27548 10382 27600
rect 23566 27548 23572 27600
rect 23624 27588 23630 27600
rect 23624 27560 26556 27588
rect 23624 27548 23630 27560
rect 5629 27523 5687 27529
rect 5629 27489 5641 27523
rect 5675 27489 5687 27523
rect 5629 27483 5687 27489
rect 9217 27523 9275 27529
rect 9217 27489 9229 27523
rect 9263 27489 9275 27523
rect 9398 27520 9404 27532
rect 9359 27492 9404 27520
rect 9217 27483 9275 27489
rect 9398 27480 9404 27492
rect 9456 27480 9462 27532
rect 9490 27480 9496 27532
rect 9548 27520 9554 27532
rect 9677 27523 9735 27529
rect 9677 27520 9689 27523
rect 9548 27492 9689 27520
rect 9548 27480 9554 27492
rect 9677 27489 9689 27492
rect 9723 27489 9735 27523
rect 9677 27483 9735 27489
rect 26053 27523 26111 27529
rect 26053 27489 26065 27523
rect 26099 27520 26111 27523
rect 26234 27520 26240 27532
rect 26099 27492 26240 27520
rect 26099 27489 26111 27492
rect 26053 27483 26111 27489
rect 26234 27480 26240 27492
rect 26292 27480 26298 27532
rect 26528 27529 26556 27560
rect 26513 27523 26571 27529
rect 26513 27489 26525 27523
rect 26559 27489 26571 27523
rect 26513 27483 26571 27489
rect 12802 27384 12808 27396
rect 12406 27356 12808 27384
rect 4062 27276 4068 27328
rect 4120 27316 4126 27328
rect 12406 27316 12434 27356
rect 12802 27344 12808 27356
rect 12860 27344 12866 27396
rect 26237 27387 26295 27393
rect 26237 27353 26249 27387
rect 26283 27384 26295 27387
rect 27062 27384 27068 27396
rect 26283 27356 27068 27384
rect 26283 27353 26295 27356
rect 26237 27347 26295 27353
rect 27062 27344 27068 27356
rect 27120 27344 27126 27396
rect 4120 27288 12434 27316
rect 4120 27276 4126 27288
rect 1104 27226 68816 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 68816 27226
rect 1104 27152 68816 27174
rect 1104 26682 68816 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 68816 26682
rect 1104 26608 68816 26630
rect 8938 26256 8944 26308
rect 8996 26296 9002 26308
rect 9490 26296 9496 26308
rect 8996 26268 9496 26296
rect 8996 26256 9002 26268
rect 9490 26256 9496 26268
rect 9548 26256 9554 26308
rect 4062 26188 4068 26240
rect 4120 26228 4126 26240
rect 23566 26228 23572 26240
rect 4120 26200 23572 26228
rect 4120 26188 4126 26200
rect 23566 26188 23572 26200
rect 23624 26188 23630 26240
rect 1104 26138 68816 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 68816 26138
rect 1104 26064 68816 26086
rect 34698 25888 34704 25900
rect 34659 25860 34704 25888
rect 34698 25848 34704 25860
rect 34756 25848 34762 25900
rect 34790 25684 34796 25696
rect 34751 25656 34796 25684
rect 34790 25644 34796 25656
rect 34848 25644 34854 25696
rect 1104 25594 68816 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 68816 25594
rect 1104 25520 68816 25542
rect 34790 25304 34796 25356
rect 34848 25344 34854 25356
rect 35069 25347 35127 25353
rect 35069 25344 35081 25347
rect 34848 25316 35081 25344
rect 34848 25304 34854 25316
rect 35069 25313 35081 25316
rect 35115 25313 35127 25347
rect 35069 25307 35127 25313
rect 34882 25276 34888 25288
rect 34843 25248 34888 25276
rect 34882 25236 34888 25248
rect 34940 25236 34946 25288
rect 36722 25208 36728 25220
rect 36683 25180 36728 25208
rect 36722 25168 36728 25180
rect 36780 25168 36786 25220
rect 1104 25050 68816 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 68816 25050
rect 1104 24976 68816 24998
rect 28810 24800 28816 24812
rect 28771 24772 28816 24800
rect 28810 24760 28816 24772
rect 28868 24760 28874 24812
rect 34882 24760 34888 24812
rect 34940 24800 34946 24812
rect 35161 24803 35219 24809
rect 35161 24800 35173 24803
rect 34940 24772 35173 24800
rect 34940 24760 34946 24772
rect 35161 24769 35173 24772
rect 35207 24769 35219 24803
rect 35161 24763 35219 24769
rect 28350 24596 28356 24608
rect 28311 24568 28356 24596
rect 28350 24556 28356 24568
rect 28408 24556 28414 24608
rect 28534 24556 28540 24608
rect 28592 24596 28598 24608
rect 28905 24599 28963 24605
rect 28905 24596 28917 24599
rect 28592 24568 28917 24596
rect 28592 24556 28598 24568
rect 28905 24565 28917 24568
rect 28951 24565 28963 24599
rect 28905 24559 28963 24565
rect 1104 24506 68816 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 68816 24506
rect 1104 24432 68816 24454
rect 58158 24148 58164 24200
rect 58216 24188 58222 24200
rect 58437 24191 58495 24197
rect 58437 24188 58449 24191
rect 58216 24160 58449 24188
rect 58216 24148 58222 24160
rect 58437 24157 58449 24160
rect 58483 24157 58495 24191
rect 58437 24151 58495 24157
rect 1104 23962 68816 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 68816 23962
rect 1104 23888 68816 23910
rect 28534 23780 28540 23792
rect 28495 23752 28540 23780
rect 28534 23740 28540 23752
rect 28592 23740 28598 23792
rect 28350 23712 28356 23724
rect 28311 23684 28356 23712
rect 28350 23672 28356 23684
rect 28408 23672 28414 23724
rect 58158 23712 58164 23724
rect 58119 23684 58164 23712
rect 58158 23672 58164 23684
rect 58216 23672 58222 23724
rect 6914 23604 6920 23656
rect 6972 23644 6978 23656
rect 28813 23647 28871 23653
rect 28813 23644 28825 23647
rect 6972 23616 28825 23644
rect 6972 23604 6978 23616
rect 28813 23613 28825 23616
rect 28859 23613 28871 23647
rect 58342 23644 58348 23656
rect 58303 23616 58348 23644
rect 28813 23607 28871 23613
rect 58342 23604 58348 23616
rect 58400 23604 58406 23656
rect 60001 23647 60059 23653
rect 60001 23613 60013 23647
rect 60047 23644 60059 23647
rect 65978 23644 65984 23656
rect 60047 23616 65984 23644
rect 60047 23613 60059 23616
rect 60001 23607 60059 23613
rect 65978 23604 65984 23616
rect 66036 23604 66042 23656
rect 1104 23418 68816 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 68816 23418
rect 1104 23344 68816 23366
rect 36722 23264 36728 23316
rect 36780 23304 36786 23316
rect 57977 23307 58035 23313
rect 36780 23276 45554 23304
rect 36780 23264 36786 23276
rect 45526 23236 45554 23276
rect 57977 23273 57989 23307
rect 58023 23304 58035 23307
rect 58342 23304 58348 23316
rect 58023 23276 58348 23304
rect 58023 23273 58035 23276
rect 57977 23267 58035 23273
rect 58342 23264 58348 23276
rect 58400 23264 58406 23316
rect 66162 23236 66168 23248
rect 45526 23208 66168 23236
rect 66162 23196 66168 23208
rect 66220 23196 66226 23248
rect 10778 23100 10784 23112
rect 10739 23072 10784 23100
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 11606 23100 11612 23112
rect 11567 23072 11612 23100
rect 11606 23060 11612 23072
rect 11664 23060 11670 23112
rect 57882 23100 57888 23112
rect 57843 23072 57888 23100
rect 57882 23060 57888 23072
rect 57940 23060 57946 23112
rect 60734 23100 60740 23112
rect 60695 23072 60740 23100
rect 60734 23060 60740 23072
rect 60792 23060 60798 23112
rect 61565 23103 61623 23109
rect 61565 23069 61577 23103
rect 61611 23069 61623 23103
rect 61565 23063 61623 23069
rect 60642 22992 60648 23044
rect 60700 23032 60706 23044
rect 61580 23032 61608 23063
rect 60700 23004 61608 23032
rect 60700 22992 60706 23004
rect 10778 22924 10784 22976
rect 10836 22964 10842 22976
rect 10873 22967 10931 22973
rect 10873 22964 10885 22967
rect 10836 22936 10885 22964
rect 10836 22924 10842 22936
rect 10873 22933 10885 22936
rect 10919 22933 10931 22967
rect 60826 22964 60832 22976
rect 60787 22936 60832 22964
rect 10873 22927 10931 22933
rect 60826 22924 60832 22936
rect 60884 22924 60890 22976
rect 1104 22874 68816 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 68816 22874
rect 1104 22800 68816 22822
rect 60826 22692 60832 22704
rect 60787 22664 60832 22692
rect 60826 22652 60832 22664
rect 60884 22652 60890 22704
rect 47578 22584 47584 22636
rect 47636 22624 47642 22636
rect 50525 22627 50583 22633
rect 50525 22624 50537 22627
rect 47636 22596 50537 22624
rect 47636 22584 47642 22596
rect 50525 22593 50537 22596
rect 50571 22624 50583 22627
rect 57882 22624 57888 22636
rect 50571 22596 57888 22624
rect 50571 22593 50583 22596
rect 50525 22587 50583 22593
rect 57882 22584 57888 22596
rect 57940 22584 57946 22636
rect 60642 22624 60648 22636
rect 60603 22596 60648 22624
rect 60642 22584 60648 22596
rect 60700 22584 60706 22636
rect 62482 22556 62488 22568
rect 62443 22528 62488 22556
rect 62482 22516 62488 22528
rect 62540 22516 62546 22568
rect 4706 22420 4712 22432
rect 4667 22392 4712 22420
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 50522 22380 50528 22432
rect 50580 22420 50586 22432
rect 50617 22423 50675 22429
rect 50617 22420 50629 22423
rect 50580 22392 50629 22420
rect 50580 22380 50586 22392
rect 50617 22389 50629 22392
rect 50663 22389 50675 22423
rect 51350 22420 51356 22432
rect 51311 22392 51356 22420
rect 50617 22383 50675 22389
rect 51350 22380 51356 22392
rect 51408 22380 51414 22432
rect 1104 22330 68816 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 68816 22330
rect 1104 22256 68816 22278
rect 3326 22108 3332 22160
rect 3384 22148 3390 22160
rect 3384 22120 5028 22148
rect 3384 22108 3390 22120
rect 4525 22083 4583 22089
rect 4525 22049 4537 22083
rect 4571 22080 4583 22083
rect 4706 22080 4712 22092
rect 4571 22052 4712 22080
rect 4571 22049 4583 22052
rect 4525 22043 4583 22049
rect 4706 22040 4712 22052
rect 4764 22040 4770 22092
rect 5000 22089 5028 22120
rect 4985 22083 5043 22089
rect 4985 22049 4997 22083
rect 5031 22049 5043 22083
rect 10778 22080 10784 22092
rect 10739 22052 10784 22080
rect 4985 22043 5043 22049
rect 10778 22040 10784 22052
rect 10836 22040 10842 22092
rect 12342 22080 12348 22092
rect 12303 22052 12348 22080
rect 12342 22040 12348 22052
rect 12400 22040 12406 22092
rect 50522 22080 50528 22092
rect 50483 22052 50528 22080
rect 50522 22040 50528 22052
rect 50580 22040 50586 22092
rect 50798 22080 50804 22092
rect 50759 22052 50804 22080
rect 50798 22040 50804 22052
rect 50856 22040 50862 22092
rect 10597 22015 10655 22021
rect 10597 21981 10609 22015
rect 10643 21981 10655 22015
rect 10597 21975 10655 21981
rect 50341 22015 50399 22021
rect 50341 21981 50353 22015
rect 50387 21981 50399 22015
rect 62942 22012 62948 22024
rect 62903 21984 62948 22012
rect 50341 21975 50399 21981
rect 4709 21947 4767 21953
rect 4709 21913 4721 21947
rect 4755 21944 4767 21947
rect 5074 21944 5080 21956
rect 4755 21916 5080 21944
rect 4755 21913 4767 21916
rect 4709 21907 4767 21913
rect 5074 21904 5080 21916
rect 5132 21904 5138 21956
rect 10612 21944 10640 21975
rect 11606 21944 11612 21956
rect 10612 21916 11612 21944
rect 11606 21904 11612 21916
rect 11664 21904 11670 21956
rect 50356 21944 50384 21975
rect 62942 21972 62948 21984
rect 63000 21972 63006 22024
rect 51350 21944 51356 21956
rect 50356 21916 51356 21944
rect 51350 21904 51356 21916
rect 51408 21904 51414 21956
rect 63037 21879 63095 21885
rect 63037 21845 63049 21879
rect 63083 21876 63095 21879
rect 63310 21876 63316 21888
rect 63083 21848 63316 21876
rect 63083 21845 63095 21848
rect 63037 21839 63095 21845
rect 63310 21836 63316 21848
rect 63368 21836 63374 21888
rect 1104 21786 68816 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 68816 21786
rect 1104 21712 68816 21734
rect 5074 21672 5080 21684
rect 5035 21644 5080 21672
rect 5074 21632 5080 21644
rect 5132 21632 5138 21684
rect 63310 21604 63316 21616
rect 63271 21576 63316 21604
rect 63310 21564 63316 21576
rect 63368 21564 63374 21616
rect 4890 21496 4896 21548
rect 4948 21536 4954 21548
rect 4985 21539 5043 21545
rect 4985 21536 4997 21539
rect 4948 21508 4997 21536
rect 4948 21496 4954 21508
rect 4985 21505 4997 21508
rect 5031 21505 5043 21539
rect 4985 21499 5043 21505
rect 63126 21468 63132 21480
rect 63087 21440 63132 21468
rect 63126 21428 63132 21440
rect 63184 21428 63190 21480
rect 64969 21471 65027 21477
rect 64969 21437 64981 21471
rect 65015 21468 65027 21471
rect 66070 21468 66076 21480
rect 65015 21440 66076 21468
rect 65015 21437 65027 21440
rect 64969 21431 65027 21437
rect 66070 21428 66076 21440
rect 66128 21428 66134 21480
rect 1104 21242 68816 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 68816 21242
rect 1104 21168 68816 21190
rect 63126 21088 63132 21140
rect 63184 21128 63190 21140
rect 63313 21131 63371 21137
rect 63313 21128 63325 21131
rect 63184 21100 63325 21128
rect 63184 21088 63190 21100
rect 63313 21097 63325 21100
rect 63359 21097 63371 21131
rect 63313 21091 63371 21097
rect 49786 20748 49792 20800
rect 49844 20788 49850 20800
rect 50798 20788 50804 20800
rect 49844 20760 50804 20788
rect 49844 20748 49850 20760
rect 50798 20748 50804 20760
rect 50856 20748 50862 20800
rect 1104 20698 68816 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 68816 20698
rect 1104 20624 68816 20646
rect 1104 20154 68816 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 68816 20154
rect 1104 20080 68816 20102
rect 32122 19796 32128 19848
rect 32180 19836 32186 19848
rect 32309 19839 32367 19845
rect 32309 19836 32321 19839
rect 32180 19808 32321 19836
rect 32180 19796 32186 19808
rect 32309 19805 32321 19808
rect 32355 19805 32367 19839
rect 32309 19799 32367 19805
rect 1104 19610 68816 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 68816 19610
rect 1104 19536 68816 19558
rect 3510 19388 3516 19440
rect 3568 19428 3574 19440
rect 33965 19431 34023 19437
rect 33965 19428 33977 19431
rect 3568 19400 33977 19428
rect 3568 19388 3574 19400
rect 33965 19397 33977 19400
rect 34011 19397 34023 19431
rect 33965 19391 34023 19397
rect 32122 19360 32128 19372
rect 32083 19332 32128 19360
rect 32122 19320 32128 19332
rect 32180 19320 32186 19372
rect 32306 19292 32312 19304
rect 32267 19264 32312 19292
rect 32306 19252 32312 19264
rect 32364 19252 32370 19304
rect 1104 19066 68816 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 68816 19066
rect 1104 18992 68816 19014
rect 32306 18912 32312 18964
rect 32364 18952 32370 18964
rect 32493 18955 32551 18961
rect 32493 18952 32505 18955
rect 32364 18924 32505 18952
rect 32364 18912 32370 18924
rect 32493 18921 32505 18924
rect 32539 18921 32551 18955
rect 32493 18915 32551 18921
rect 32401 18751 32459 18757
rect 32401 18717 32413 18751
rect 32447 18748 32459 18751
rect 45370 18748 45376 18760
rect 32447 18720 45376 18748
rect 32447 18717 32459 18720
rect 32401 18711 32459 18717
rect 45370 18708 45376 18720
rect 45428 18708 45434 18760
rect 1104 18522 68816 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 68816 18522
rect 1104 18448 68816 18470
rect 5442 18068 5448 18080
rect 5403 18040 5448 18068
rect 5442 18028 5448 18040
rect 5500 18028 5506 18080
rect 1104 17978 68816 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 68816 17978
rect 1104 17904 68816 17926
rect 5169 17731 5227 17737
rect 5169 17697 5181 17731
rect 5215 17728 5227 17731
rect 5442 17728 5448 17740
rect 5215 17700 5448 17728
rect 5215 17697 5227 17700
rect 5169 17691 5227 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 6822 17728 6828 17740
rect 6783 17700 6828 17728
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 62669 17663 62727 17669
rect 62669 17629 62681 17663
rect 62715 17660 62727 17663
rect 62942 17660 62948 17672
rect 62715 17632 62948 17660
rect 62715 17629 62727 17632
rect 62669 17623 62727 17629
rect 62942 17620 62948 17632
rect 63000 17620 63006 17672
rect 63034 17620 63040 17672
rect 63092 17660 63098 17672
rect 63497 17663 63555 17669
rect 63497 17660 63509 17663
rect 63092 17632 63509 17660
rect 63092 17620 63098 17632
rect 63497 17629 63509 17632
rect 63543 17629 63555 17663
rect 63497 17623 63555 17629
rect 5353 17595 5411 17601
rect 5353 17561 5365 17595
rect 5399 17592 5411 17595
rect 5534 17592 5540 17604
rect 5399 17564 5540 17592
rect 5399 17561 5411 17564
rect 5353 17555 5411 17561
rect 5534 17552 5540 17564
rect 5592 17552 5598 17604
rect 62761 17527 62819 17533
rect 62761 17493 62773 17527
rect 62807 17524 62819 17527
rect 63218 17524 63224 17536
rect 62807 17496 63224 17524
rect 62807 17493 62819 17496
rect 62761 17487 62819 17493
rect 63218 17484 63224 17496
rect 63276 17484 63282 17536
rect 1104 17434 68816 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 68816 17434
rect 1104 17360 68816 17382
rect 5534 17320 5540 17332
rect 5495 17292 5540 17320
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 63218 17252 63224 17264
rect 63179 17224 63224 17252
rect 63218 17212 63224 17224
rect 63276 17212 63282 17264
rect 4890 17144 4896 17196
rect 4948 17184 4954 17196
rect 5442 17184 5448 17196
rect 4948 17156 5448 17184
rect 4948 17144 4954 17156
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 63034 17184 63040 17196
rect 62995 17156 63040 17184
rect 63034 17144 63040 17156
rect 63092 17144 63098 17196
rect 64782 17116 64788 17128
rect 64743 17088 64788 17116
rect 64782 17076 64788 17088
rect 64840 17076 64846 17128
rect 1104 16890 68816 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 68816 16890
rect 1104 16816 68816 16838
rect 3326 16532 3332 16584
rect 3384 16572 3390 16584
rect 8938 16572 8944 16584
rect 3384 16544 8944 16572
rect 3384 16532 3390 16544
rect 8938 16532 8944 16544
rect 8996 16532 9002 16584
rect 1104 16346 68816 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 68816 16346
rect 1104 16272 68816 16294
rect 1104 15802 68816 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 68816 15802
rect 1104 15728 68816 15750
rect 12802 15444 12808 15496
rect 12860 15484 12866 15496
rect 13081 15487 13139 15493
rect 13081 15484 13093 15487
rect 12860 15456 13093 15484
rect 12860 15444 12866 15456
rect 13081 15453 13093 15456
rect 13127 15453 13139 15487
rect 13081 15447 13139 15453
rect 1104 15258 68816 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 68816 15258
rect 1104 15184 68816 15206
rect 62482 15104 62488 15156
rect 62540 15144 62546 15156
rect 66070 15144 66076 15156
rect 62540 15116 66076 15144
rect 62540 15104 62546 15116
rect 66070 15104 66076 15116
rect 66128 15104 66134 15156
rect 12802 15008 12808 15020
rect 12763 14980 12808 15008
rect 12802 14968 12808 14980
rect 12860 14968 12866 15020
rect 12986 14940 12992 14952
rect 12947 14912 12992 14940
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 13538 14940 13544 14952
rect 13499 14912 13544 14940
rect 13538 14900 13544 14912
rect 13596 14900 13602 14952
rect 1104 14714 68816 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 68816 14714
rect 1104 14640 68816 14662
rect 12897 14603 12955 14609
rect 12897 14569 12909 14603
rect 12943 14600 12955 14603
rect 12986 14600 12992 14612
rect 12943 14572 12992 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 5442 14356 5448 14408
rect 5500 14396 5506 14408
rect 12805 14399 12863 14405
rect 12805 14396 12817 14399
rect 5500 14368 12817 14396
rect 5500 14356 5506 14368
rect 12805 14365 12817 14368
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 19426 14356 19432 14408
rect 19484 14396 19490 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 19484 14368 19625 14396
rect 19484 14356 19490 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 22094 14396 22100 14408
rect 22055 14368 22100 14396
rect 19613 14359 19671 14365
rect 22094 14356 22100 14368
rect 22152 14356 22158 14408
rect 22186 14260 22192 14272
rect 22147 14232 22192 14260
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 1104 14170 68816 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 68816 14170
rect 1104 14096 68816 14118
rect 22186 13988 22192 14000
rect 22147 13960 22192 13988
rect 22186 13948 22192 13960
rect 22244 13948 22250 14000
rect 19426 13920 19432 13932
rect 19387 13892 19432 13920
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 19610 13852 19616 13864
rect 19571 13824 19616 13852
rect 19610 13812 19616 13824
rect 19668 13812 19674 13864
rect 19889 13855 19947 13861
rect 19889 13852 19901 13855
rect 19720 13824 19901 13852
rect 3326 13744 3332 13796
rect 3384 13784 3390 13796
rect 19720 13784 19748 13824
rect 19889 13821 19901 13824
rect 19935 13821 19947 13855
rect 19889 13815 19947 13821
rect 22005 13855 22063 13861
rect 22005 13821 22017 13855
rect 22051 13852 22063 13855
rect 22186 13852 22192 13864
rect 22051 13824 22192 13852
rect 22051 13821 22063 13824
rect 22005 13815 22063 13821
rect 22186 13812 22192 13824
rect 22244 13812 22250 13864
rect 22554 13852 22560 13864
rect 22515 13824 22560 13852
rect 22554 13812 22560 13824
rect 22612 13812 22618 13864
rect 3384 13756 19748 13784
rect 3384 13744 3390 13756
rect 1104 13626 68816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 68816 13626
rect 1104 13552 68816 13574
rect 19610 13472 19616 13524
rect 19668 13512 19674 13524
rect 19981 13515 20039 13521
rect 19981 13512 19993 13515
rect 19668 13484 19993 13512
rect 19668 13472 19674 13484
rect 19981 13481 19993 13484
rect 20027 13481 20039 13515
rect 22186 13512 22192 13524
rect 22147 13484 22192 13512
rect 19981 13475 20039 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13308 19947 13311
rect 22094 13308 22100 13320
rect 19935 13280 22100 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 22094 13268 22100 13280
rect 22152 13308 22158 13320
rect 35529 13311 35587 13317
rect 35529 13308 35541 13311
rect 22152 13280 35541 13308
rect 22152 13268 22158 13280
rect 35529 13277 35541 13280
rect 35575 13277 35587 13311
rect 35529 13271 35587 13277
rect 35618 13172 35624 13184
rect 35579 13144 35624 13172
rect 35618 13132 35624 13144
rect 35676 13132 35682 13184
rect 1104 13082 68816 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 68816 13082
rect 1104 13008 68816 13030
rect 35434 12588 35440 12640
rect 35492 12628 35498 12640
rect 35713 12631 35771 12637
rect 35713 12628 35725 12631
rect 35492 12600 35725 12628
rect 35492 12588 35498 12600
rect 35713 12597 35725 12600
rect 35759 12597 35771 12631
rect 35713 12591 35771 12597
rect 1104 12538 68816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 68816 12538
rect 1104 12464 68816 12486
rect 45278 12356 45284 12368
rect 34808 12328 45284 12356
rect 26878 12180 26884 12232
rect 26936 12220 26942 12232
rect 34701 12223 34759 12229
rect 34701 12220 34713 12223
rect 26936 12192 34713 12220
rect 26936 12180 26942 12192
rect 34701 12189 34713 12192
rect 34747 12220 34759 12223
rect 34808 12220 34836 12328
rect 45278 12316 45284 12328
rect 45336 12316 45342 12368
rect 35434 12288 35440 12300
rect 35395 12260 35440 12288
rect 35434 12248 35440 12260
rect 35492 12248 35498 12300
rect 35618 12288 35624 12300
rect 35579 12260 35624 12288
rect 35618 12248 35624 12260
rect 35676 12248 35682 12300
rect 36078 12288 36084 12300
rect 36039 12260 36084 12288
rect 36078 12248 36084 12260
rect 36136 12248 36142 12300
rect 34747 12192 34836 12220
rect 34747 12189 34759 12192
rect 34701 12183 34759 12189
rect 63402 12180 63408 12232
rect 63460 12220 63466 12232
rect 63589 12223 63647 12229
rect 63589 12220 63601 12223
rect 63460 12192 63601 12220
rect 63460 12180 63466 12192
rect 63589 12189 63601 12192
rect 63635 12189 63647 12223
rect 63589 12183 63647 12189
rect 34422 12044 34428 12096
rect 34480 12084 34486 12096
rect 34793 12087 34851 12093
rect 34793 12084 34805 12087
rect 34480 12056 34805 12084
rect 34480 12044 34486 12056
rect 34793 12053 34805 12056
rect 34839 12053 34851 12087
rect 34793 12047 34851 12053
rect 1104 11994 68816 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 68816 11994
rect 1104 11920 68816 11942
rect 34422 11812 34428 11824
rect 34383 11784 34428 11812
rect 34422 11772 34428 11784
rect 34480 11772 34486 11824
rect 63402 11744 63408 11756
rect 63363 11716 63408 11744
rect 63402 11704 63408 11716
rect 63460 11704 63466 11756
rect 33781 11679 33839 11685
rect 33781 11645 33793 11679
rect 33827 11676 33839 11679
rect 34241 11679 34299 11685
rect 34241 11676 34253 11679
rect 33827 11648 34253 11676
rect 33827 11645 33839 11648
rect 33781 11639 33839 11645
rect 34241 11645 34253 11648
rect 34287 11645 34299 11679
rect 34790 11676 34796 11688
rect 34751 11648 34796 11676
rect 34241 11639 34299 11645
rect 34790 11636 34796 11648
rect 34848 11636 34854 11688
rect 63310 11636 63316 11688
rect 63368 11676 63374 11688
rect 63589 11679 63647 11685
rect 63589 11676 63601 11679
rect 63368 11648 63601 11676
rect 63368 11636 63374 11648
rect 63589 11645 63601 11648
rect 63635 11645 63647 11679
rect 65242 11676 65248 11688
rect 65203 11648 65248 11676
rect 63589 11639 63647 11645
rect 65242 11636 65248 11648
rect 65300 11636 65306 11688
rect 24578 11500 24584 11552
rect 24636 11540 24642 11552
rect 24765 11543 24823 11549
rect 24765 11540 24777 11543
rect 24636 11512 24777 11540
rect 24636 11500 24642 11512
rect 24765 11509 24777 11512
rect 24811 11509 24823 11543
rect 24765 11503 24823 11509
rect 30098 11500 30104 11552
rect 30156 11540 30162 11552
rect 30285 11543 30343 11549
rect 30285 11540 30297 11543
rect 30156 11512 30297 11540
rect 30156 11500 30162 11512
rect 30285 11509 30297 11512
rect 30331 11509 30343 11543
rect 30285 11503 30343 11509
rect 1104 11450 68816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 68816 11450
rect 1104 11376 68816 11398
rect 63310 11336 63316 11348
rect 63271 11308 63316 11336
rect 63310 11296 63316 11308
rect 63368 11296 63374 11348
rect 5810 11228 5816 11280
rect 5868 11268 5874 11280
rect 5868 11240 35388 11268
rect 5868 11228 5874 11240
rect 3602 11160 3608 11212
rect 3660 11200 3666 11212
rect 35360 11209 35388 11240
rect 30561 11203 30619 11209
rect 30561 11200 30573 11203
rect 3660 11172 30573 11200
rect 3660 11160 3666 11172
rect 30561 11169 30573 11172
rect 30607 11169 30619 11203
rect 30561 11163 30619 11169
rect 35345 11203 35403 11209
rect 35345 11169 35357 11203
rect 35391 11169 35403 11203
rect 35345 11163 35403 11169
rect 24578 11132 24584 11144
rect 24539 11104 24584 11132
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 26878 11132 26884 11144
rect 26839 11104 26884 11132
rect 26878 11092 26884 11104
rect 26936 11092 26942 11144
rect 30098 11132 30104 11144
rect 30059 11104 30104 11132
rect 30098 11092 30104 11104
rect 30156 11092 30162 11144
rect 34149 11135 34207 11141
rect 34149 11101 34161 11135
rect 34195 11132 34207 11135
rect 34885 11135 34943 11141
rect 34885 11132 34897 11135
rect 34195 11104 34897 11132
rect 34195 11101 34207 11104
rect 34149 11095 34207 11101
rect 34885 11101 34897 11104
rect 34931 11101 34943 11135
rect 34885 11095 34943 11101
rect 63221 11135 63279 11141
rect 63221 11101 63233 11135
rect 63267 11132 63279 11135
rect 63678 11132 63684 11144
rect 63267 11104 63684 11132
rect 63267 11101 63279 11104
rect 63221 11095 63279 11101
rect 63678 11092 63684 11104
rect 63736 11092 63742 11144
rect 19978 11024 19984 11076
rect 20036 11064 20042 11076
rect 20036 11036 24716 11064
rect 20036 11024 20042 11036
rect 24688 10996 24716 11036
rect 24762 11024 24768 11076
rect 24820 11064 24826 11076
rect 26421 11067 26479 11073
rect 26421 11064 26433 11067
rect 24820 11036 24865 11064
rect 24964 11036 26433 11064
rect 24820 11024 24826 11036
rect 24964 10996 24992 11036
rect 26421 11033 26433 11036
rect 26467 11033 26479 11067
rect 26421 11027 26479 11033
rect 30285 11067 30343 11073
rect 30285 11033 30297 11067
rect 30331 11064 30343 11067
rect 30650 11064 30656 11076
rect 30331 11036 30656 11064
rect 30331 11033 30343 11036
rect 30285 11027 30343 11033
rect 30650 11024 30656 11036
rect 30708 11024 30714 11076
rect 35066 11064 35072 11076
rect 35027 11036 35072 11064
rect 35066 11024 35072 11036
rect 35124 11024 35130 11076
rect 24688 10968 24992 10996
rect 26234 10956 26240 11008
rect 26292 10996 26298 11008
rect 26973 10999 27031 11005
rect 26973 10996 26985 10999
rect 26292 10968 26985 10996
rect 26292 10956 26298 10968
rect 26973 10965 26985 10968
rect 27019 10965 27031 10999
rect 26973 10959 27031 10965
rect 1104 10906 68816 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 68816 10906
rect 1104 10832 68816 10854
rect 24854 10752 24860 10804
rect 24912 10792 24918 10804
rect 25133 10795 25191 10801
rect 25133 10792 25145 10795
rect 24912 10764 25145 10792
rect 24912 10752 24918 10764
rect 25133 10761 25145 10764
rect 25179 10761 25191 10795
rect 30650 10792 30656 10804
rect 30611 10764 30656 10792
rect 25133 10755 25191 10761
rect 30650 10752 30656 10764
rect 30708 10752 30714 10804
rect 35066 10752 35072 10804
rect 35124 10792 35130 10804
rect 35253 10795 35311 10801
rect 35253 10792 35265 10795
rect 35124 10764 35265 10792
rect 35124 10752 35130 10764
rect 35253 10761 35265 10764
rect 35299 10761 35311 10795
rect 35253 10755 35311 10761
rect 25041 10659 25099 10665
rect 25041 10625 25053 10659
rect 25087 10656 25099 10659
rect 26878 10656 26884 10668
rect 25087 10628 26884 10656
rect 25087 10625 25099 10628
rect 25041 10619 25099 10625
rect 26878 10616 26884 10628
rect 26936 10616 26942 10668
rect 30561 10659 30619 10665
rect 30561 10625 30573 10659
rect 30607 10656 30619 10659
rect 35161 10659 35219 10665
rect 35161 10656 35173 10659
rect 30607 10628 35173 10656
rect 30607 10625 30619 10628
rect 30561 10619 30619 10625
rect 35161 10625 35173 10628
rect 35207 10656 35219 10659
rect 48958 10656 48964 10668
rect 35207 10628 48964 10656
rect 35207 10625 35219 10628
rect 35161 10619 35219 10625
rect 48958 10616 48964 10628
rect 49016 10616 49022 10668
rect 26050 10412 26056 10464
rect 26108 10452 26114 10464
rect 26329 10455 26387 10461
rect 26329 10452 26341 10455
rect 26108 10424 26341 10452
rect 26108 10412 26114 10424
rect 26329 10421 26341 10424
rect 26375 10421 26387 10455
rect 26329 10415 26387 10421
rect 1104 10362 68816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 68816 10362
rect 1104 10288 68816 10310
rect 26050 10112 26056 10124
rect 26011 10084 26056 10112
rect 26050 10072 26056 10084
rect 26108 10072 26114 10124
rect 26234 10112 26240 10124
rect 26195 10084 26240 10112
rect 26234 10072 26240 10084
rect 26292 10072 26298 10124
rect 43346 10044 43352 10056
rect 43307 10016 43352 10044
rect 43346 10004 43352 10016
rect 43404 10044 43410 10056
rect 54386 10044 54392 10056
rect 43404 10016 54392 10044
rect 43404 10004 43410 10016
rect 54386 10004 54392 10016
rect 54444 10004 54450 10056
rect 27798 9936 27804 9988
rect 27856 9976 27862 9988
rect 27893 9979 27951 9985
rect 27893 9976 27905 9979
rect 27856 9948 27905 9976
rect 27856 9936 27862 9948
rect 27893 9945 27905 9948
rect 27939 9945 27951 9979
rect 27893 9939 27951 9945
rect 43438 9908 43444 9920
rect 43399 9880 43444 9908
rect 43438 9868 43444 9880
rect 43496 9868 43502 9920
rect 1104 9818 68816 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 68816 9818
rect 1104 9744 68816 9766
rect 43438 9636 43444 9648
rect 43399 9608 43444 9636
rect 43438 9596 43444 9608
rect 43496 9596 43502 9648
rect 43257 9503 43315 9509
rect 43257 9469 43269 9503
rect 43303 9500 43315 9503
rect 43530 9500 43536 9512
rect 43303 9472 43536 9500
rect 43303 9469 43315 9472
rect 43257 9463 43315 9469
rect 43530 9460 43536 9472
rect 43588 9460 43594 9512
rect 43806 9500 43812 9512
rect 43767 9472 43812 9500
rect 43806 9460 43812 9472
rect 43864 9460 43870 9512
rect 1104 9274 68816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 68816 9274
rect 1104 9200 68816 9222
rect 43530 9160 43536 9172
rect 43491 9132 43536 9160
rect 43530 9120 43536 9132
rect 43588 9120 43594 9172
rect 26881 9027 26939 9033
rect 26881 9024 26893 9027
rect 6886 8996 26893 9024
rect 14 8848 20 8900
rect 72 8888 78 8900
rect 6886 8888 6914 8996
rect 26881 8993 26893 8996
rect 26927 8993 26939 9027
rect 26881 8987 26939 8993
rect 25961 8959 26019 8965
rect 25961 8925 25973 8959
rect 26007 8956 26019 8959
rect 26421 8959 26479 8965
rect 26421 8956 26433 8959
rect 26007 8928 26433 8956
rect 26007 8925 26019 8928
rect 25961 8919 26019 8925
rect 26421 8925 26433 8928
rect 26467 8925 26479 8959
rect 54386 8956 54392 8968
rect 54347 8928 54392 8956
rect 26421 8919 26479 8925
rect 54386 8916 54392 8928
rect 54444 8916 54450 8968
rect 54754 8916 54760 8968
rect 54812 8956 54818 8968
rect 55493 8959 55551 8965
rect 55493 8956 55505 8959
rect 54812 8928 55505 8956
rect 54812 8916 54818 8928
rect 55493 8925 55505 8928
rect 55539 8925 55551 8959
rect 55493 8919 55551 8925
rect 72 8860 6914 8888
rect 26605 8891 26663 8897
rect 72 8848 78 8860
rect 26605 8857 26617 8891
rect 26651 8888 26663 8891
rect 27062 8888 27068 8900
rect 26651 8860 27068 8888
rect 26651 8857 26663 8860
rect 26605 8851 26663 8857
rect 27062 8848 27068 8860
rect 27120 8848 27126 8900
rect 54481 8823 54539 8829
rect 54481 8789 54493 8823
rect 54527 8820 54539 8823
rect 54938 8820 54944 8832
rect 54527 8792 54944 8820
rect 54527 8789 54539 8792
rect 54481 8783 54539 8789
rect 54938 8780 54944 8792
rect 54996 8780 55002 8832
rect 1104 8730 68816 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 68816 8730
rect 1104 8656 68816 8678
rect 27062 8616 27068 8628
rect 27023 8588 27068 8616
rect 27062 8576 27068 8588
rect 27120 8576 27126 8628
rect 54938 8548 54944 8560
rect 54899 8520 54944 8548
rect 54938 8508 54944 8520
rect 54996 8508 55002 8560
rect 26973 8483 27031 8489
rect 26973 8449 26985 8483
rect 27019 8480 27031 8483
rect 43346 8480 43352 8492
rect 27019 8452 43352 8480
rect 27019 8449 27031 8452
rect 26973 8443 27031 8449
rect 43346 8440 43352 8452
rect 43404 8440 43410 8492
rect 54754 8480 54760 8492
rect 54715 8452 54760 8480
rect 54754 8440 54760 8452
rect 54812 8440 54818 8492
rect 56597 8415 56655 8421
rect 56597 8381 56609 8415
rect 56643 8412 56655 8415
rect 59262 8412 59268 8424
rect 56643 8384 59268 8412
rect 56643 8381 56655 8384
rect 56597 8375 56655 8381
rect 59262 8372 59268 8384
rect 59320 8372 59326 8424
rect 1104 8186 68816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 68816 8186
rect 1104 8112 68816 8134
rect 1104 7642 68816 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 68816 7642
rect 1104 7568 68816 7590
rect 1104 7098 68816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 68816 7098
rect 1104 7024 68816 7046
rect 1104 6554 68816 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 68816 6554
rect 1104 6480 68816 6502
rect 1104 6010 68816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 68816 6010
rect 1104 5936 68816 5958
rect 1104 5466 68816 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 68816 5466
rect 1104 5392 68816 5414
rect 1104 4922 68816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 68816 4922
rect 1104 4848 68816 4870
rect 1104 4378 68816 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 68816 4378
rect 1104 4304 68816 4326
rect 45186 4088 45192 4140
rect 45244 4128 45250 4140
rect 47026 4128 47032 4140
rect 45244 4100 47032 4128
rect 45244 4088 45250 4100
rect 47026 4088 47032 4100
rect 47084 4088 47090 4140
rect 45094 4020 45100 4072
rect 45152 4060 45158 4072
rect 46842 4060 46848 4072
rect 45152 4032 46848 4060
rect 45152 4020 45158 4032
rect 46842 4020 46848 4032
rect 46900 4020 46906 4072
rect 1104 3834 68816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 68816 3834
rect 1104 3760 68816 3782
rect 24486 3544 24492 3596
rect 24544 3584 24550 3596
rect 27341 3587 27399 3593
rect 27341 3584 27353 3587
rect 24544 3556 27353 3584
rect 24544 3544 24550 3556
rect 27341 3553 27353 3556
rect 27387 3553 27399 3587
rect 27341 3547 27399 3553
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 68922 3584 68928 3596
rect 28960 3556 68928 3584
rect 28960 3544 28966 3556
rect 68922 3544 68928 3556
rect 68980 3544 68986 3596
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 6822 3516 6828 3528
rect 4672 3488 6828 3516
rect 4672 3476 4678 3488
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 12342 3516 12348 3528
rect 11020 3488 12348 3516
rect 11020 3476 11026 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 26418 3476 26424 3528
rect 26476 3516 26482 3528
rect 26881 3519 26939 3525
rect 26881 3516 26893 3519
rect 26476 3488 26893 3516
rect 26476 3476 26482 3488
rect 26881 3485 26893 3488
rect 26927 3485 26939 3519
rect 40678 3516 40684 3528
rect 40639 3488 40684 3516
rect 26881 3479 26939 3485
rect 40678 3476 40684 3488
rect 40736 3476 40742 3528
rect 67818 3476 67824 3528
rect 67876 3516 67882 3528
rect 69566 3516 69572 3528
rect 67876 3488 69572 3516
rect 67876 3476 67882 3488
rect 69566 3476 69572 3488
rect 69624 3476 69630 3528
rect 27062 3448 27068 3460
rect 27023 3420 27068 3448
rect 27062 3408 27068 3420
rect 27120 3408 27126 3460
rect 40865 3451 40923 3457
rect 40865 3417 40877 3451
rect 40911 3448 40923 3451
rect 41782 3448 41788 3460
rect 40911 3420 41788 3448
rect 40911 3417 40923 3420
rect 40865 3411 40923 3417
rect 41782 3408 41788 3420
rect 41840 3408 41846 3460
rect 42521 3451 42579 3457
rect 42521 3417 42533 3451
rect 42567 3417 42579 3451
rect 42521 3411 42579 3417
rect 41230 3340 41236 3392
rect 41288 3380 41294 3392
rect 42536 3380 42564 3411
rect 45462 3408 45468 3460
rect 45520 3448 45526 3460
rect 61194 3448 61200 3460
rect 45520 3420 61200 3448
rect 45520 3408 45526 3420
rect 61194 3408 61200 3420
rect 61252 3408 61258 3460
rect 41288 3352 42564 3380
rect 41288 3340 41294 3352
rect 1104 3290 68816 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 68816 3290
rect 1104 3216 68816 3238
rect 41782 3176 41788 3188
rect 41743 3148 41788 3176
rect 41782 3136 41788 3148
rect 41840 3136 41846 3188
rect 56502 3136 56508 3188
rect 56560 3176 56566 3188
rect 62482 3176 62488 3188
rect 56560 3148 62488 3176
rect 56560 3136 56566 3148
rect 62482 3136 62488 3148
rect 62540 3136 62546 3188
rect 27065 3111 27123 3117
rect 27065 3077 27077 3111
rect 27111 3108 27123 3111
rect 27801 3111 27859 3117
rect 27801 3108 27813 3111
rect 27111 3080 27813 3108
rect 27111 3077 27123 3080
rect 27065 3071 27123 3077
rect 27801 3077 27813 3080
rect 27847 3077 27859 3111
rect 27801 3071 27859 3077
rect 26418 3040 26424 3052
rect 26379 3012 26424 3040
rect 26418 3000 26424 3012
rect 26476 3000 26482 3052
rect 26970 3040 26976 3052
rect 26931 3012 26976 3040
rect 26970 3000 26976 3012
rect 27028 3000 27034 3052
rect 41690 3040 41696 3052
rect 41603 3012 41696 3040
rect 41690 3000 41696 3012
rect 41748 3040 41754 3052
rect 42978 3040 42984 3052
rect 41748 3012 42984 3040
rect 41748 3000 41754 3012
rect 42978 3000 42984 3012
rect 43036 3000 43042 3052
rect 27614 2972 27620 2984
rect 27575 2944 27620 2972
rect 27614 2932 27620 2944
rect 27672 2932 27678 2984
rect 28077 2975 28135 2981
rect 28077 2941 28089 2975
rect 28123 2941 28135 2975
rect 28077 2935 28135 2941
rect 38933 2975 38991 2981
rect 38933 2941 38945 2975
rect 38979 2972 38991 2975
rect 39393 2975 39451 2981
rect 39393 2972 39405 2975
rect 38979 2944 39405 2972
rect 38979 2941 38991 2944
rect 38933 2935 38991 2941
rect 39393 2941 39405 2944
rect 39439 2941 39451 2975
rect 39574 2972 39580 2984
rect 39535 2944 39580 2972
rect 39393 2935 39451 2941
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 28092 2904 28120 2935
rect 39574 2932 39580 2944
rect 39632 2932 39638 2984
rect 39942 2972 39948 2984
rect 39903 2944 39948 2972
rect 39942 2932 39948 2944
rect 40000 2932 40006 2984
rect 14884 2876 28120 2904
rect 14884 2864 14890 2876
rect 1104 2746 68816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 68816 2746
rect 1104 2672 68816 2694
rect 27062 2592 27068 2644
rect 27120 2632 27126 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 27120 2604 27169 2632
rect 27120 2592 27126 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 27157 2595 27215 2601
rect 27614 2592 27620 2644
rect 27672 2632 27678 2644
rect 27893 2635 27951 2641
rect 27893 2632 27905 2635
rect 27672 2604 27905 2632
rect 27672 2592 27678 2604
rect 27893 2601 27905 2604
rect 27939 2601 27951 2635
rect 27893 2595 27951 2601
rect 39574 2592 39580 2644
rect 39632 2632 39638 2644
rect 39945 2635 40003 2641
rect 39945 2632 39957 2635
rect 39632 2604 39957 2632
rect 39632 2592 39638 2604
rect 39945 2601 39957 2604
rect 39991 2601 40003 2635
rect 39945 2595 40003 2601
rect 40678 2592 40684 2644
rect 40736 2632 40742 2644
rect 40865 2635 40923 2641
rect 40865 2632 40877 2635
rect 40736 2604 40877 2632
rect 40736 2592 40742 2604
rect 40865 2601 40877 2604
rect 40911 2601 40923 2635
rect 40865 2595 40923 2601
rect 26970 2388 26976 2440
rect 27028 2428 27034 2440
rect 27065 2431 27123 2437
rect 27065 2428 27077 2431
rect 27028 2400 27077 2428
rect 27028 2388 27034 2400
rect 27065 2397 27077 2400
rect 27111 2428 27123 2431
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 27111 2400 39865 2428
rect 27111 2397 27123 2400
rect 27065 2391 27123 2397
rect 39853 2397 39865 2400
rect 39899 2428 39911 2431
rect 41690 2428 41696 2440
rect 39899 2400 41696 2428
rect 39899 2397 39911 2400
rect 39853 2391 39911 2397
rect 41690 2388 41696 2400
rect 41748 2388 41754 2440
rect 1104 2202 68816 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 68816 2202
rect 1104 2128 68816 2150
rect 3418 1300 3424 1352
rect 3476 1340 3482 1352
rect 27798 1340 27804 1352
rect 3476 1312 27804 1340
rect 3476 1300 3482 1312
rect 27798 1300 27804 1312
rect 27856 1300 27862 1352
rect 59262 1300 59268 1352
rect 59320 1340 59326 1352
rect 66162 1340 66168 1352
rect 59320 1312 66168 1340
rect 59320 1300 59326 1312
rect 66162 1300 66168 1312
rect 66220 1300 66226 1352
<< via1 >>
rect 47400 71408 47452 71460
rect 48228 71408 48280 71460
rect 19574 69606 19626 69658
rect 19638 69606 19690 69658
rect 19702 69606 19754 69658
rect 19766 69606 19818 69658
rect 19830 69606 19882 69658
rect 50294 69606 50346 69658
rect 50358 69606 50410 69658
rect 50422 69606 50474 69658
rect 50486 69606 50538 69658
rect 50550 69606 50602 69658
rect 67456 69479 67508 69488
rect 67456 69445 67465 69479
rect 67465 69445 67499 69479
rect 67499 69445 67508 69479
rect 67456 69436 67508 69445
rect 1492 69411 1544 69420
rect 1492 69377 1501 69411
rect 1501 69377 1535 69411
rect 1535 69377 1544 69411
rect 1492 69368 1544 69377
rect 55404 69368 55456 69420
rect 31392 69300 31444 69352
rect 34060 69300 34112 69352
rect 30472 69232 30524 69284
rect 46756 69207 46808 69216
rect 46756 69173 46765 69207
rect 46765 69173 46799 69207
rect 46799 69173 46808 69207
rect 46756 69164 46808 69173
rect 51264 69207 51316 69216
rect 51264 69173 51273 69207
rect 51273 69173 51307 69207
rect 51307 69173 51316 69207
rect 51264 69164 51316 69173
rect 56968 69207 57020 69216
rect 56968 69173 56977 69207
rect 56977 69173 57011 69207
rect 57011 69173 57020 69207
rect 56968 69164 57020 69173
rect 58992 69164 59044 69216
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 34934 69062 34986 69114
rect 34998 69062 35050 69114
rect 35062 69062 35114 69114
rect 35126 69062 35178 69114
rect 35190 69062 35242 69114
rect 65654 69062 65706 69114
rect 65718 69062 65770 69114
rect 65782 69062 65834 69114
rect 65846 69062 65898 69114
rect 65910 69062 65962 69114
rect 25136 68960 25188 69012
rect 28264 68960 28316 69012
rect 46572 68960 46624 69012
rect 52828 68960 52880 69012
rect 64144 68960 64196 69012
rect 66996 68960 67048 69012
rect 41880 68892 41932 68944
rect 46756 68824 46808 68876
rect 56692 68892 56744 68944
rect 51264 68824 51316 68876
rect 51540 68867 51592 68876
rect 51540 68833 51549 68867
rect 51549 68833 51583 68867
rect 51583 68833 51592 68867
rect 51540 68824 51592 68833
rect 56968 68824 57020 68876
rect 49148 68756 49200 68808
rect 58900 68799 58952 68808
rect 58900 68765 58909 68799
rect 58909 68765 58943 68799
rect 58943 68765 58952 68799
rect 58900 68756 58952 68765
rect 51172 68731 51224 68740
rect 40684 68620 40736 68672
rect 46572 68620 46624 68672
rect 51172 68697 51181 68731
rect 51181 68697 51215 68731
rect 51215 68697 51224 68731
rect 51172 68688 51224 68697
rect 56416 68731 56468 68740
rect 56416 68697 56425 68731
rect 56425 68697 56459 68731
rect 56459 68697 56468 68731
rect 56416 68688 56468 68697
rect 53288 68620 53340 68672
rect 63132 68688 63184 68740
rect 59176 68620 59228 68672
rect 19574 68518 19626 68570
rect 19638 68518 19690 68570
rect 19702 68518 19754 68570
rect 19766 68518 19818 68570
rect 19830 68518 19882 68570
rect 50294 68518 50346 68570
rect 50358 68518 50410 68570
rect 50422 68518 50474 68570
rect 50486 68518 50538 68570
rect 50550 68518 50602 68570
rect 16764 68416 16816 68468
rect 33140 68416 33192 68468
rect 38568 68416 38620 68468
rect 51172 68459 51224 68468
rect 6460 68348 6512 68400
rect 22744 68348 22796 68400
rect 24124 68348 24176 68400
rect 44456 68348 44508 68400
rect 51172 68425 51181 68459
rect 51181 68425 51215 68459
rect 51215 68425 51224 68459
rect 51172 68416 51224 68425
rect 54116 68416 54168 68468
rect 56416 68459 56468 68468
rect 56416 68425 56425 68459
rect 56425 68425 56459 68459
rect 56459 68425 56468 68459
rect 56416 68416 56468 68425
rect 53380 68348 53432 68400
rect 65340 68348 65392 68400
rect 23204 68280 23256 68332
rect 29644 68280 29696 68332
rect 49148 68280 49200 68332
rect 58992 68323 59044 68332
rect 58992 68289 59001 68323
rect 59001 68289 59035 68323
rect 59035 68289 59044 68323
rect 58992 68280 59044 68289
rect 58900 68212 58952 68264
rect 59176 68255 59228 68264
rect 59176 68221 59185 68255
rect 59185 68221 59219 68255
rect 59219 68221 59228 68255
rect 59176 68212 59228 68221
rect 68284 68212 68336 68264
rect 3884 68076 3936 68128
rect 5540 68076 5592 68128
rect 30288 68076 30340 68128
rect 31116 68076 31168 68128
rect 37924 68076 37976 68128
rect 39304 68076 39356 68128
rect 58624 68076 58676 68128
rect 60556 68076 60608 68128
rect 67732 68076 67784 68128
rect 69204 68076 69256 68128
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 34934 67974 34986 68026
rect 34998 67974 35050 68026
rect 35062 67974 35114 68026
rect 35126 67974 35178 68026
rect 35190 67974 35242 68026
rect 65654 67974 65706 68026
rect 65718 67974 65770 68026
rect 65782 67974 65834 68026
rect 65846 67974 65898 68026
rect 65910 67974 65962 68026
rect 60924 67711 60976 67720
rect 60924 67677 60933 67711
rect 60933 67677 60967 67711
rect 60967 67677 60976 67711
rect 60924 67668 60976 67677
rect 43168 67600 43220 67652
rect 44180 67600 44232 67652
rect 61108 67643 61160 67652
rect 61108 67609 61117 67643
rect 61117 67609 61151 67643
rect 61151 67609 61160 67643
rect 61108 67600 61160 67609
rect 62764 67643 62816 67652
rect 62764 67609 62773 67643
rect 62773 67609 62807 67643
rect 62807 67609 62816 67643
rect 62764 67600 62816 67609
rect 19574 67430 19626 67482
rect 19638 67430 19690 67482
rect 19702 67430 19754 67482
rect 19766 67430 19818 67482
rect 19830 67430 19882 67482
rect 50294 67430 50346 67482
rect 50358 67430 50410 67482
rect 50422 67430 50474 67482
rect 50486 67430 50538 67482
rect 50550 67430 50602 67482
rect 61108 67328 61160 67380
rect 58900 67192 58952 67244
rect 60924 67192 60976 67244
rect 62764 66988 62816 67040
rect 66168 66988 66220 67040
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 37464 66580 37516 66632
rect 43812 66580 43864 66632
rect 19574 66342 19626 66394
rect 19638 66342 19690 66394
rect 19702 66342 19754 66394
rect 19766 66342 19818 66394
rect 19830 66342 19882 66394
rect 50294 66342 50346 66394
rect 50358 66342 50410 66394
rect 50422 66342 50474 66394
rect 50486 66342 50538 66394
rect 50550 66342 50602 66394
rect 37464 66147 37516 66156
rect 37464 66113 37473 66147
rect 37473 66113 37507 66147
rect 37507 66113 37516 66147
rect 37464 66104 37516 66113
rect 43812 66147 43864 66156
rect 43812 66113 43821 66147
rect 43821 66113 43855 66147
rect 43855 66113 43864 66147
rect 43812 66104 43864 66113
rect 37740 66036 37792 66088
rect 38660 66079 38712 66088
rect 38660 66045 38669 66079
rect 38669 66045 38703 66079
rect 38703 66045 38712 66079
rect 38660 66036 38712 66045
rect 43996 66079 44048 66088
rect 43996 66045 44005 66079
rect 44005 66045 44039 66079
rect 44039 66045 44048 66079
rect 43996 66036 44048 66045
rect 45468 66079 45520 66088
rect 45468 66045 45477 66079
rect 45477 66045 45511 66079
rect 45511 66045 45520 66079
rect 45468 66036 45520 66045
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 37740 65739 37792 65748
rect 37740 65705 37749 65739
rect 37749 65705 37783 65739
rect 37783 65705 37792 65739
rect 37740 65696 37792 65705
rect 43996 65696 44048 65748
rect 31392 65560 31444 65612
rect 6736 65492 6788 65544
rect 31852 65535 31904 65544
rect 31852 65501 31861 65535
rect 31861 65501 31895 65535
rect 31895 65501 31904 65535
rect 31852 65492 31904 65501
rect 42616 65492 42668 65544
rect 43904 65492 43956 65544
rect 43536 65424 43588 65476
rect 19574 65254 19626 65306
rect 19638 65254 19690 65306
rect 19702 65254 19754 65306
rect 19766 65254 19818 65306
rect 19830 65254 19882 65306
rect 50294 65254 50346 65306
rect 50358 65254 50410 65306
rect 50422 65254 50474 65306
rect 50486 65254 50538 65306
rect 50550 65254 50602 65306
rect 30932 65084 30984 65136
rect 6736 65059 6788 65068
rect 6736 65025 6745 65059
rect 6745 65025 6779 65059
rect 6779 65025 6788 65059
rect 6736 65016 6788 65025
rect 31392 65059 31444 65068
rect 31392 65025 31401 65059
rect 31401 65025 31435 65059
rect 31435 65025 31444 65059
rect 31392 65016 31444 65025
rect 42616 65059 42668 65068
rect 42616 65025 42625 65059
rect 42625 65025 42659 65059
rect 42659 65025 42668 65059
rect 42616 65016 42668 65025
rect 6920 64991 6972 65000
rect 6920 64957 6929 64991
rect 6929 64957 6963 64991
rect 6963 64957 6972 64991
rect 6920 64948 6972 64957
rect 33140 64991 33192 65000
rect 5540 64880 5592 64932
rect 33140 64957 33149 64991
rect 33149 64957 33183 64991
rect 33183 64957 33192 64991
rect 33140 64948 33192 64957
rect 42800 64991 42852 65000
rect 42800 64957 42809 64991
rect 42809 64957 42843 64991
rect 42843 64957 42852 64991
rect 42800 64948 42852 64957
rect 44180 64991 44232 65000
rect 44180 64957 44189 64991
rect 44189 64957 44223 64991
rect 44223 64957 44232 64991
rect 44180 64948 44232 64957
rect 55956 64855 56008 64864
rect 55956 64821 55965 64855
rect 55965 64821 55999 64855
rect 55999 64821 56008 64855
rect 55956 64812 56008 64821
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 34934 64710 34986 64762
rect 34998 64710 35050 64762
rect 35062 64710 35114 64762
rect 35126 64710 35178 64762
rect 35190 64710 35242 64762
rect 65654 64710 65706 64762
rect 65718 64710 65770 64762
rect 65782 64710 65834 64762
rect 65846 64710 65898 64762
rect 65910 64710 65962 64762
rect 6920 64608 6972 64660
rect 30472 64651 30524 64660
rect 30472 64617 30481 64651
rect 30481 64617 30515 64651
rect 30515 64617 30524 64651
rect 30472 64608 30524 64617
rect 30932 64651 30984 64660
rect 30932 64617 30941 64651
rect 30941 64617 30975 64651
rect 30975 64617 30984 64651
rect 30932 64608 30984 64617
rect 42800 64651 42852 64660
rect 42800 64617 42809 64651
rect 42809 64617 42843 64651
rect 42843 64617 42852 64651
rect 42800 64608 42852 64617
rect 31208 64583 31260 64592
rect 31208 64549 31217 64583
rect 31217 64549 31251 64583
rect 31251 64549 31260 64583
rect 31208 64540 31260 64549
rect 4620 64472 4672 64524
rect 31852 64472 31904 64524
rect 55956 64472 56008 64524
rect 64144 64472 64196 64524
rect 7196 64404 7248 64456
rect 29736 64447 29788 64456
rect 29736 64413 29745 64447
rect 29745 64413 29779 64447
rect 29779 64413 29788 64447
rect 29736 64404 29788 64413
rect 31576 64404 31628 64456
rect 34060 64404 34112 64456
rect 34152 64447 34204 64456
rect 34152 64413 34161 64447
rect 34161 64413 34195 64447
rect 34195 64413 34204 64447
rect 34152 64404 34204 64413
rect 43904 64404 43956 64456
rect 30840 64379 30892 64388
rect 30840 64345 30849 64379
rect 30849 64345 30883 64379
rect 30883 64345 30892 64379
rect 30840 64336 30892 64345
rect 33232 64336 33284 64388
rect 55864 64379 55916 64388
rect 55864 64345 55873 64379
rect 55873 64345 55907 64379
rect 55907 64345 55916 64379
rect 55864 64336 55916 64345
rect 19574 64166 19626 64218
rect 19638 64166 19690 64218
rect 19702 64166 19754 64218
rect 19766 64166 19818 64218
rect 19830 64166 19882 64218
rect 50294 64166 50346 64218
rect 50358 64166 50410 64218
rect 50422 64166 50474 64218
rect 50486 64166 50538 64218
rect 50550 64166 50602 64218
rect 30840 64064 30892 64116
rect 32588 64064 32640 64116
rect 55864 64064 55916 64116
rect 31116 64039 31168 64048
rect 31116 64005 31125 64039
rect 31125 64005 31159 64039
rect 31159 64005 31168 64039
rect 31116 63996 31168 64005
rect 37924 63996 37976 64048
rect 31576 63928 31628 63980
rect 55588 63971 55640 63980
rect 55588 63937 55597 63971
rect 55597 63937 55631 63971
rect 55631 63937 55640 63971
rect 55588 63928 55640 63937
rect 28724 63860 28776 63912
rect 29736 63860 29788 63912
rect 32312 63903 32364 63912
rect 32312 63869 32321 63903
rect 32321 63869 32355 63903
rect 32355 63869 32364 63903
rect 32312 63860 32364 63869
rect 58072 63767 58124 63776
rect 58072 63733 58081 63767
rect 58081 63733 58115 63767
rect 58115 63733 58124 63767
rect 58072 63724 58124 63733
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 34934 63622 34986 63674
rect 34998 63622 35050 63674
rect 35062 63622 35114 63674
rect 35126 63622 35178 63674
rect 35190 63622 35242 63674
rect 65654 63622 65706 63674
rect 65718 63622 65770 63674
rect 65782 63622 65834 63674
rect 65846 63622 65898 63674
rect 65910 63622 65962 63674
rect 28724 63520 28776 63572
rect 30656 63520 30708 63572
rect 33232 63495 33284 63504
rect 33232 63461 33241 63495
rect 33241 63461 33275 63495
rect 33275 63461 33284 63495
rect 33232 63452 33284 63461
rect 29644 63384 29696 63436
rect 58072 63384 58124 63436
rect 59084 63427 59136 63436
rect 59084 63393 59093 63427
rect 59093 63393 59127 63427
rect 59127 63393 59136 63427
rect 59084 63384 59136 63393
rect 30656 63359 30708 63368
rect 30656 63325 30665 63359
rect 30665 63325 30699 63359
rect 30699 63325 30708 63359
rect 30656 63316 30708 63325
rect 31208 63316 31260 63368
rect 33140 63359 33192 63368
rect 33140 63325 33149 63359
rect 33149 63325 33183 63359
rect 33183 63325 33192 63359
rect 33140 63316 33192 63325
rect 44180 63316 44232 63368
rect 49700 63316 49752 63368
rect 32312 63248 32364 63300
rect 57980 63248 58032 63300
rect 32588 63180 32640 63232
rect 19574 63078 19626 63130
rect 19638 63078 19690 63130
rect 19702 63078 19754 63130
rect 19766 63078 19818 63130
rect 19830 63078 19882 63130
rect 50294 63078 50346 63130
rect 50358 63078 50410 63130
rect 50422 63078 50474 63130
rect 50486 63078 50538 63130
rect 50550 63078 50602 63130
rect 49148 63019 49200 63028
rect 49148 62985 49157 63019
rect 49157 62985 49191 63019
rect 49191 62985 49200 63019
rect 49148 62976 49200 62985
rect 57980 63019 58032 63028
rect 57980 62985 57989 63019
rect 57989 62985 58023 63019
rect 58023 62985 58032 63019
rect 57980 62976 58032 62985
rect 49516 62840 49568 62892
rect 49700 62883 49752 62892
rect 49700 62849 49709 62883
rect 49709 62849 49743 62883
rect 49743 62849 49752 62883
rect 49700 62840 49752 62849
rect 64512 62840 64564 62892
rect 32404 62772 32456 62824
rect 30564 62704 30616 62756
rect 50252 62772 50304 62824
rect 49792 62704 49844 62756
rect 65156 62704 65208 62756
rect 46480 62636 46532 62688
rect 65340 62636 65392 62688
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 34934 62534 34986 62586
rect 34998 62534 35050 62586
rect 35062 62534 35114 62586
rect 35126 62534 35178 62586
rect 35190 62534 35242 62586
rect 65654 62534 65706 62586
rect 65718 62534 65770 62586
rect 65782 62534 65834 62586
rect 65846 62534 65898 62586
rect 65910 62534 65962 62586
rect 32404 62475 32456 62484
rect 32404 62441 32413 62475
rect 32413 62441 32447 62475
rect 32447 62441 32456 62475
rect 32404 62432 32456 62441
rect 50252 62475 50304 62484
rect 50252 62441 50261 62475
rect 50261 62441 50295 62475
rect 50295 62441 50304 62475
rect 50252 62432 50304 62441
rect 46480 62339 46532 62348
rect 46480 62305 46489 62339
rect 46489 62305 46523 62339
rect 46523 62305 46532 62339
rect 46480 62296 46532 62305
rect 48228 62339 48280 62348
rect 48228 62305 48237 62339
rect 48237 62305 48271 62339
rect 48271 62305 48280 62339
rect 48228 62296 48280 62305
rect 67456 62339 67508 62348
rect 67456 62305 67465 62339
rect 67465 62305 67499 62339
rect 67499 62305 67508 62339
rect 67456 62296 67508 62305
rect 33140 62228 33192 62280
rect 46664 62203 46716 62212
rect 46664 62169 46673 62203
rect 46673 62169 46707 62203
rect 46707 62169 46716 62203
rect 46664 62160 46716 62169
rect 38476 62092 38528 62144
rect 54484 62228 54536 62280
rect 65800 62203 65852 62212
rect 65800 62169 65809 62203
rect 65809 62169 65843 62203
rect 65843 62169 65852 62203
rect 65800 62160 65852 62169
rect 19574 61990 19626 62042
rect 19638 61990 19690 62042
rect 19702 61990 19754 62042
rect 19766 61990 19818 62042
rect 19830 61990 19882 62042
rect 50294 61990 50346 62042
rect 50358 61990 50410 62042
rect 50422 61990 50474 62042
rect 50486 61990 50538 62042
rect 50550 61990 50602 62042
rect 46664 61931 46716 61940
rect 46664 61897 46673 61931
rect 46673 61897 46707 61931
rect 46707 61897 46716 61931
rect 46664 61888 46716 61897
rect 65800 61888 65852 61940
rect 37280 61752 37332 61804
rect 55588 61820 55640 61872
rect 65340 61863 65392 61872
rect 65340 61829 65349 61863
rect 65349 61829 65383 61863
rect 65383 61829 65392 61863
rect 65340 61820 65392 61829
rect 67732 61820 67784 61872
rect 54484 61795 54536 61804
rect 54484 61761 54493 61795
rect 54493 61761 54527 61795
rect 54527 61761 54536 61795
rect 54484 61752 54536 61761
rect 64512 61795 64564 61804
rect 64512 61761 64521 61795
rect 64521 61761 64555 61795
rect 64555 61761 64564 61795
rect 64512 61752 64564 61761
rect 65156 61795 65208 61804
rect 65156 61761 65165 61795
rect 65165 61761 65199 61795
rect 65199 61761 65208 61795
rect 65156 61752 65208 61761
rect 54668 61727 54720 61736
rect 54668 61693 54677 61727
rect 54677 61693 54711 61727
rect 54711 61693 54720 61727
rect 54668 61684 54720 61693
rect 66076 61684 66128 61736
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 65654 61446 65706 61498
rect 65718 61446 65770 61498
rect 65782 61446 65834 61498
rect 65846 61446 65898 61498
rect 65910 61446 65962 61498
rect 54668 61344 54720 61396
rect 23020 61140 23072 61192
rect 44180 61140 44232 61192
rect 44364 61140 44416 61192
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 23020 60707 23072 60716
rect 23020 60673 23029 60707
rect 23029 60673 23063 60707
rect 23063 60673 23072 60707
rect 23020 60664 23072 60673
rect 1400 60639 1452 60648
rect 1400 60605 1409 60639
rect 1409 60605 1443 60639
rect 1443 60605 1452 60639
rect 1400 60596 1452 60605
rect 23572 60596 23624 60648
rect 23664 60639 23716 60648
rect 23664 60605 23673 60639
rect 23673 60605 23707 60639
rect 23707 60605 23716 60639
rect 23664 60596 23716 60605
rect 34152 60528 34204 60580
rect 22744 60460 22796 60512
rect 23388 60460 23440 60512
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 65654 60358 65706 60410
rect 65718 60358 65770 60410
rect 65782 60358 65834 60410
rect 65846 60358 65898 60410
rect 65910 60358 65962 60410
rect 23572 60299 23624 60308
rect 23572 60265 23581 60299
rect 23581 60265 23615 60299
rect 23615 60265 23624 60299
rect 23572 60256 23624 60265
rect 47216 60188 47268 60240
rect 24860 60052 24912 60104
rect 26976 60095 27028 60104
rect 26976 60061 26985 60095
rect 26985 60061 27019 60095
rect 27019 60061 27028 60095
rect 26976 60052 27028 60061
rect 47676 59984 47728 60036
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 47676 59755 47728 59764
rect 47676 59721 47685 59755
rect 47685 59721 47719 59755
rect 47719 59721 47728 59755
rect 47676 59712 47728 59721
rect 28816 59687 28868 59696
rect 28816 59653 28825 59687
rect 28825 59653 28859 59687
rect 28859 59653 28868 59687
rect 28816 59644 28868 59653
rect 48504 59576 48556 59628
rect 27160 59551 27212 59560
rect 27160 59517 27169 59551
rect 27169 59517 27203 59551
rect 27203 59517 27212 59551
rect 27160 59508 27212 59517
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 65654 59270 65706 59322
rect 65718 59270 65770 59322
rect 65782 59270 65834 59322
rect 65846 59270 65898 59322
rect 65910 59270 65962 59322
rect 27160 59168 27212 59220
rect 3332 58896 3384 58948
rect 26976 59032 27028 59084
rect 24952 58964 25004 59016
rect 27160 58896 27212 58948
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 27160 58667 27212 58676
rect 27160 58633 27169 58667
rect 27169 58633 27203 58667
rect 27203 58633 27212 58667
rect 27160 58624 27212 58633
rect 24860 58488 24912 58540
rect 37924 58488 37976 58540
rect 38476 58488 38528 58540
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 65654 58182 65706 58234
rect 65718 58182 65770 58234
rect 65782 58182 65834 58234
rect 65846 58182 65898 58234
rect 65910 58182 65962 58234
rect 48412 57876 48464 57928
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 48412 57443 48464 57452
rect 48412 57409 48421 57443
rect 48421 57409 48455 57443
rect 48455 57409 48464 57443
rect 48412 57400 48464 57409
rect 48596 57375 48648 57384
rect 48596 57341 48605 57375
rect 48605 57341 48639 57375
rect 48639 57341 48648 57375
rect 48596 57332 48648 57341
rect 48320 57264 48372 57316
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 48596 57035 48648 57044
rect 48596 57001 48605 57035
rect 48605 57001 48639 57035
rect 48639 57001 48648 57035
rect 48596 56992 48648 57001
rect 11060 56856 11112 56908
rect 48504 56831 48556 56840
rect 48504 56797 48513 56831
rect 48513 56797 48547 56831
rect 48547 56797 48556 56831
rect 48504 56788 48556 56797
rect 49056 56788 49108 56840
rect 11336 56763 11388 56772
rect 11336 56729 11345 56763
rect 11345 56729 11379 56763
rect 11379 56729 11388 56763
rect 11336 56720 11388 56729
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 11336 56448 11388 56500
rect 20628 56448 20680 56500
rect 24952 56448 25004 56500
rect 11520 56355 11572 56364
rect 11520 56321 11529 56355
rect 11529 56321 11563 56355
rect 11563 56321 11572 56355
rect 11520 56312 11572 56321
rect 20628 56312 20680 56364
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 57888 55700 57940 55752
rect 2964 55564 3016 55616
rect 33048 55564 33100 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 32588 55267 32640 55276
rect 32588 55233 32597 55267
rect 32597 55233 32631 55267
rect 32631 55233 32640 55267
rect 32588 55224 32640 55233
rect 37280 55267 37332 55276
rect 37280 55233 37289 55267
rect 37289 55233 37323 55267
rect 37323 55233 37332 55267
rect 37280 55224 37332 55233
rect 49056 55224 49108 55276
rect 57888 55267 57940 55276
rect 57888 55233 57897 55267
rect 57897 55233 57931 55267
rect 57931 55233 57940 55267
rect 57888 55224 57940 55233
rect 33048 55199 33100 55208
rect 33048 55165 33057 55199
rect 33057 55165 33091 55199
rect 33091 55165 33100 55199
rect 33048 55156 33100 55165
rect 66076 55156 66128 55208
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 2780 54000 2832 54052
rect 5724 54000 5776 54052
rect 27528 53975 27580 53984
rect 27528 53941 27537 53975
rect 27537 53941 27571 53975
rect 27571 53941 27580 53975
rect 27528 53932 27580 53941
rect 38844 53932 38896 53984
rect 51448 53975 51500 53984
rect 51448 53941 51457 53975
rect 51457 53941 51491 53975
rect 51491 53941 51500 53975
rect 51448 53932 51500 53941
rect 66260 53932 66312 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 3516 53592 3568 53644
rect 27528 53592 27580 53644
rect 66168 53660 66220 53712
rect 51448 53592 51500 53644
rect 66260 53635 66312 53644
rect 66260 53601 66269 53635
rect 66269 53601 66303 53635
rect 66303 53601 66312 53635
rect 66260 53592 66312 53601
rect 27896 53456 27948 53508
rect 51356 53499 51408 53508
rect 51356 53465 51365 53499
rect 51365 53465 51399 53499
rect 51399 53465 51408 53499
rect 51356 53456 51408 53465
rect 58624 53456 58676 53508
rect 66444 53499 66496 53508
rect 66444 53465 66453 53499
rect 66453 53465 66487 53499
rect 66487 53465 66496 53499
rect 66444 53456 66496 53465
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 27896 53227 27948 53236
rect 27896 53193 27905 53227
rect 27905 53193 27939 53227
rect 27939 53193 27948 53227
rect 27896 53184 27948 53193
rect 51356 53184 51408 53236
rect 66444 53184 66496 53236
rect 40684 53159 40736 53168
rect 40684 53125 40693 53159
rect 40693 53125 40727 53159
rect 40727 53125 40736 53159
rect 40684 53116 40736 53125
rect 38200 53091 38252 53100
rect 38200 53057 38209 53091
rect 38209 53057 38243 53091
rect 38243 53057 38252 53091
rect 38200 53048 38252 53057
rect 38844 53091 38896 53100
rect 38844 53057 38853 53091
rect 38853 53057 38887 53091
rect 38887 53057 38896 53091
rect 38844 53048 38896 53057
rect 51080 53091 51132 53100
rect 51080 53057 51089 53091
rect 51089 53057 51123 53091
rect 51123 53057 51132 53091
rect 51080 53048 51132 53057
rect 67456 53091 67508 53100
rect 67456 53057 67465 53091
rect 67465 53057 67499 53091
rect 67499 53057 67508 53091
rect 67456 53048 67508 53057
rect 45376 52912 45428 52964
rect 5264 52844 5316 52896
rect 7564 52844 7616 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 5264 52547 5316 52556
rect 5264 52513 5273 52547
rect 5273 52513 5307 52547
rect 5307 52513 5316 52547
rect 5264 52504 5316 52513
rect 5632 52504 5684 52556
rect 5724 52547 5776 52556
rect 5724 52513 5733 52547
rect 5733 52513 5767 52547
rect 5767 52513 5776 52547
rect 5724 52504 5776 52513
rect 11520 52436 11572 52488
rect 7748 52300 7800 52352
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 5632 52096 5684 52148
rect 2964 52028 3016 52080
rect 7748 52071 7800 52080
rect 7748 52037 7757 52071
rect 7757 52037 7791 52071
rect 7791 52037 7800 52071
rect 7748 52028 7800 52037
rect 7564 52003 7616 52012
rect 7564 51969 7573 52003
rect 7573 51969 7607 52003
rect 7607 51969 7616 52003
rect 7564 51960 7616 51969
rect 20904 51824 20956 51876
rect 51356 51756 51408 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 51356 51459 51408 51468
rect 51356 51425 51365 51459
rect 51365 51425 51399 51459
rect 51399 51425 51408 51459
rect 51356 51416 51408 51425
rect 53288 51416 53340 51468
rect 34888 51348 34940 51400
rect 45560 51391 45612 51400
rect 45560 51357 45569 51391
rect 45569 51357 45603 51391
rect 45603 51357 45612 51391
rect 45560 51348 45612 51357
rect 51540 51323 51592 51332
rect 51540 51289 51549 51323
rect 51549 51289 51583 51323
rect 51583 51289 51592 51323
rect 51540 51280 51592 51289
rect 36728 51212 36780 51264
rect 66076 51212 66128 51264
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 51540 51008 51592 51060
rect 3332 50940 3384 50992
rect 36728 50983 36780 50992
rect 34888 50915 34940 50924
rect 34888 50881 34897 50915
rect 34897 50881 34931 50915
rect 34931 50881 34940 50915
rect 34888 50872 34940 50881
rect 35348 50804 35400 50856
rect 36728 50949 36737 50983
rect 36737 50949 36771 50983
rect 36771 50949 36780 50983
rect 36728 50940 36780 50949
rect 45560 50940 45612 50992
rect 53196 50872 53248 50924
rect 45560 50804 45612 50856
rect 63224 50668 63276 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 35348 50507 35400 50516
rect 35348 50473 35357 50507
rect 35357 50473 35391 50507
rect 35391 50473 35400 50507
rect 35348 50464 35400 50473
rect 45560 50464 45612 50516
rect 63224 50371 63276 50380
rect 63224 50337 63233 50371
rect 63233 50337 63267 50371
rect 63267 50337 63276 50371
rect 63224 50328 63276 50337
rect 64788 50371 64840 50380
rect 64788 50337 64797 50371
rect 64797 50337 64831 50371
rect 64831 50337 64840 50371
rect 64788 50328 64840 50337
rect 6920 50260 6972 50312
rect 27436 50260 27488 50312
rect 29736 50260 29788 50312
rect 35440 50260 35492 50312
rect 38200 50260 38252 50312
rect 47584 50260 47636 50312
rect 63408 50235 63460 50244
rect 63408 50201 63417 50235
rect 63417 50201 63451 50235
rect 63451 50201 63460 50235
rect 63408 50192 63460 50201
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 28264 49920 28316 49972
rect 29276 49895 29328 49904
rect 29276 49861 29285 49895
rect 29285 49861 29319 49895
rect 29319 49861 29328 49895
rect 29276 49852 29328 49861
rect 63408 49920 63460 49972
rect 6920 49827 6972 49836
rect 6920 49793 6929 49827
rect 6929 49793 6963 49827
rect 6963 49793 6972 49827
rect 6920 49784 6972 49793
rect 27436 49827 27488 49836
rect 27436 49793 27445 49827
rect 27445 49793 27479 49827
rect 27479 49793 27488 49827
rect 27436 49784 27488 49793
rect 29736 49827 29788 49836
rect 29736 49793 29745 49827
rect 29745 49793 29779 49827
rect 29779 49793 29788 49827
rect 29736 49784 29788 49793
rect 4068 49716 4120 49768
rect 7104 49759 7156 49768
rect 7104 49725 7113 49759
rect 7113 49725 7147 49759
rect 7147 49725 7156 49759
rect 7104 49716 7156 49725
rect 27620 49759 27672 49768
rect 27620 49725 27629 49759
rect 27629 49725 27663 49759
rect 27663 49725 27672 49759
rect 27620 49716 27672 49725
rect 30380 49716 30432 49768
rect 62948 49784 63000 49836
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 7104 49376 7156 49428
rect 27620 49376 27672 49428
rect 30380 49419 30432 49428
rect 30380 49385 30389 49419
rect 30389 49385 30423 49419
rect 30423 49385 30432 49419
rect 30380 49376 30432 49385
rect 7196 49215 7248 49224
rect 7196 49181 7205 49215
rect 7205 49181 7239 49215
rect 7239 49181 7248 49215
rect 7196 49172 7248 49181
rect 28540 49215 28592 49224
rect 28540 49181 28549 49215
rect 28549 49181 28583 49215
rect 28583 49181 28592 49215
rect 28540 49172 28592 49181
rect 41604 49172 41656 49224
rect 53840 49172 53892 49224
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 44364 48764 44416 48816
rect 64696 48764 64748 48816
rect 44180 48739 44232 48748
rect 44180 48705 44189 48739
rect 44189 48705 44223 48739
rect 44223 48705 44232 48739
rect 44180 48696 44232 48705
rect 53196 48739 53248 48748
rect 53196 48705 53205 48739
rect 53205 48705 53239 48739
rect 53239 48705 53248 48739
rect 53196 48696 53248 48705
rect 53840 48739 53892 48748
rect 53840 48705 53849 48739
rect 53849 48705 53883 48739
rect 53883 48705 53892 48739
rect 53840 48696 53892 48705
rect 64512 48560 64564 48612
rect 64696 48560 64748 48612
rect 43628 48535 43680 48544
rect 43628 48501 43637 48535
rect 43637 48501 43671 48535
rect 43671 48501 43680 48535
rect 43628 48492 43680 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 43904 48220 43956 48272
rect 43444 48084 43496 48136
rect 44180 48016 44232 48068
rect 45284 48059 45336 48068
rect 45284 48025 45293 48059
rect 45293 48025 45327 48059
rect 45327 48025 45336 48059
rect 45284 48016 45336 48025
rect 53196 48016 53248 48068
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 43628 47719 43680 47728
rect 43628 47685 43637 47719
rect 43637 47685 43671 47719
rect 43671 47685 43680 47719
rect 43628 47676 43680 47685
rect 43444 47651 43496 47660
rect 43444 47617 43453 47651
rect 43453 47617 43487 47651
rect 43487 47617 43496 47651
rect 43444 47608 43496 47617
rect 64696 47651 64748 47660
rect 64696 47617 64705 47651
rect 64705 47617 64739 47651
rect 64739 47617 64748 47651
rect 64696 47608 64748 47617
rect 4068 47540 4120 47592
rect 65340 47583 65392 47592
rect 65340 47549 65349 47583
rect 65349 47549 65383 47583
rect 65383 47549 65392 47583
rect 65340 47540 65392 47549
rect 67180 47583 67232 47592
rect 67180 47549 67189 47583
rect 67189 47549 67223 47583
rect 67223 47549 67232 47583
rect 67180 47540 67232 47549
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 65340 47200 65392 47252
rect 43536 47064 43588 47116
rect 43812 47064 43864 47116
rect 44180 47064 44232 47116
rect 45376 47107 45428 47116
rect 45376 47073 45385 47107
rect 45385 47073 45419 47107
rect 45419 47073 45428 47107
rect 45376 47064 45428 47073
rect 62948 46928 63000 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 37280 45908 37332 45960
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 37280 45475 37332 45484
rect 37280 45441 37289 45475
rect 37289 45441 37323 45475
rect 37323 45441 37332 45475
rect 37280 45432 37332 45441
rect 48780 45432 48832 45484
rect 49516 45475 49568 45484
rect 49516 45441 49525 45475
rect 49525 45441 49559 45475
rect 49559 45441 49568 45475
rect 49516 45432 49568 45441
rect 37464 45407 37516 45416
rect 37464 45373 37473 45407
rect 37473 45373 37507 45407
rect 37507 45373 37516 45407
rect 37464 45364 37516 45373
rect 38476 45407 38528 45416
rect 38476 45373 38485 45407
rect 38485 45373 38519 45407
rect 38519 45373 38528 45407
rect 38476 45364 38528 45373
rect 47584 45296 47636 45348
rect 67456 45296 67508 45348
rect 14740 45228 14792 45280
rect 66260 45228 66312 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 37464 45024 37516 45076
rect 3424 44956 3476 45008
rect 14740 44931 14792 44940
rect 14740 44897 14749 44931
rect 14749 44897 14783 44931
rect 14783 44897 14792 44931
rect 14740 44888 14792 44897
rect 66260 44931 66312 44940
rect 66260 44897 66269 44931
rect 66269 44897 66303 44931
rect 66303 44897 66312 44931
rect 66260 44888 66312 44897
rect 68100 44931 68152 44940
rect 68100 44897 68109 44931
rect 68109 44897 68143 44931
rect 68143 44897 68152 44931
rect 68100 44888 68152 44897
rect 22192 44820 22244 44872
rect 28540 44820 28592 44872
rect 15108 44752 15160 44804
rect 66444 44795 66496 44804
rect 66444 44761 66453 44795
rect 66453 44761 66487 44795
rect 66487 44761 66496 44795
rect 66444 44752 66496 44761
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 15108 44523 15160 44532
rect 15108 44489 15117 44523
rect 15117 44489 15151 44523
rect 15151 44489 15160 44523
rect 15108 44480 15160 44489
rect 66444 44480 66496 44532
rect 13728 44344 13780 44396
rect 37740 44387 37792 44396
rect 37740 44353 37749 44387
rect 37749 44353 37783 44387
rect 37783 44353 37792 44387
rect 37740 44344 37792 44353
rect 43812 44344 43864 44396
rect 67456 44387 67508 44396
rect 67456 44353 67465 44387
rect 67465 44353 67499 44387
rect 67499 44353 67508 44387
rect 67456 44344 67508 44353
rect 37924 44276 37976 44328
rect 52092 44276 52144 44328
rect 44088 44140 44140 44192
rect 48780 44140 48832 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 52092 43775 52144 43784
rect 52092 43741 52101 43775
rect 52101 43741 52135 43775
rect 52135 43741 52144 43775
rect 52092 43732 52144 43741
rect 52736 43775 52788 43784
rect 52736 43741 52745 43775
rect 52745 43741 52779 43775
rect 52779 43741 52788 43775
rect 52736 43732 52788 43741
rect 66168 43664 66220 43716
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 52736 43256 52788 43308
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 52092 42644 52144 42696
rect 54944 42508 54996 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 54944 42279 54996 42288
rect 54944 42245 54953 42279
rect 54953 42245 54987 42279
rect 54987 42245 54996 42279
rect 54944 42236 54996 42245
rect 12624 42168 12676 42220
rect 13728 42168 13780 42220
rect 44088 42211 44140 42220
rect 20628 42100 20680 42152
rect 24860 42100 24912 42152
rect 44088 42177 44097 42211
rect 44097 42177 44131 42211
rect 44131 42177 44140 42211
rect 44088 42168 44140 42177
rect 37740 42100 37792 42152
rect 43536 42100 43588 42152
rect 56508 42143 56560 42152
rect 56508 42109 56517 42143
rect 56517 42109 56551 42143
rect 56551 42109 56560 42143
rect 56508 42100 56560 42109
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 24860 41420 24912 41472
rect 26424 41420 26476 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 44364 41080 44416 41132
rect 57888 41055 57940 41064
rect 57888 41021 57897 41055
rect 57897 41021 57931 41055
rect 57931 41021 57940 41055
rect 57888 41012 57940 41021
rect 66168 41012 66220 41064
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 57888 40715 57940 40724
rect 57888 40681 57897 40715
rect 57897 40681 57931 40715
rect 57931 40681 57940 40715
rect 57888 40672 57940 40681
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 3056 40060 3108 40112
rect 23848 40060 23900 40112
rect 9588 39788 9640 39840
rect 35348 39831 35400 39840
rect 35348 39797 35357 39831
rect 35357 39797 35391 39831
rect 35391 39797 35400 39831
rect 35348 39788 35400 39797
rect 60464 39788 60516 39840
rect 63224 39788 63276 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 3332 39312 3384 39364
rect 9588 39491 9640 39500
rect 9588 39457 9597 39491
rect 9597 39457 9631 39491
rect 9631 39457 9640 39491
rect 9588 39448 9640 39457
rect 22100 39448 22152 39500
rect 35348 39448 35400 39500
rect 36912 39491 36964 39500
rect 36912 39457 36921 39491
rect 36921 39457 36955 39491
rect 36955 39457 36964 39491
rect 36912 39448 36964 39457
rect 60464 39491 60516 39500
rect 60464 39457 60473 39491
rect 60473 39457 60507 39491
rect 60507 39457 60516 39491
rect 60464 39448 60516 39457
rect 62028 39491 62080 39500
rect 62028 39457 62037 39491
rect 62037 39457 62071 39491
rect 62071 39457 62080 39491
rect 62028 39448 62080 39457
rect 63224 39491 63276 39500
rect 63224 39457 63233 39491
rect 63233 39457 63267 39491
rect 63267 39457 63276 39491
rect 63224 39448 63276 39457
rect 64788 39491 64840 39500
rect 64788 39457 64797 39491
rect 64797 39457 64831 39491
rect 64831 39457 64840 39491
rect 64788 39448 64840 39457
rect 22284 39380 22336 39432
rect 9864 39312 9916 39364
rect 34888 39312 34940 39364
rect 60648 39355 60700 39364
rect 60648 39321 60657 39355
rect 60657 39321 60691 39355
rect 60691 39321 60700 39355
rect 60648 39312 60700 39321
rect 63500 39312 63552 39364
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 9864 39083 9916 39092
rect 9864 39049 9873 39083
rect 9873 39049 9907 39083
rect 9907 39049 9916 39083
rect 9864 39040 9916 39049
rect 34888 39083 34940 39092
rect 34888 39049 34897 39083
rect 34897 39049 34931 39083
rect 34931 39049 34940 39083
rect 34888 39040 34940 39049
rect 60648 39040 60700 39092
rect 63500 39083 63552 39092
rect 63500 39049 63509 39083
rect 63509 39049 63543 39083
rect 63543 39049 63552 39083
rect 63500 39040 63552 39049
rect 24124 39015 24176 39024
rect 24124 38981 24133 39015
rect 24133 38981 24167 39015
rect 24167 38981 24176 39015
rect 24124 38972 24176 38981
rect 9772 38947 9824 38956
rect 9772 38913 9781 38947
rect 9781 38913 9815 38947
rect 9815 38913 9824 38947
rect 9772 38904 9824 38913
rect 22284 38947 22336 38956
rect 22284 38913 22293 38947
rect 22293 38913 22327 38947
rect 22327 38913 22336 38947
rect 22284 38904 22336 38913
rect 34704 38904 34756 38956
rect 44364 38904 44416 38956
rect 48780 38972 48832 39024
rect 22468 38879 22520 38888
rect 22468 38845 22477 38879
rect 22477 38845 22511 38879
rect 22511 38845 22520 38879
rect 22468 38836 22520 38845
rect 46388 38836 46440 38888
rect 61844 38904 61896 38956
rect 63408 38947 63460 38956
rect 63408 38913 63417 38947
rect 63417 38913 63451 38947
rect 63451 38913 63460 38947
rect 63408 38904 63460 38913
rect 45192 38700 45244 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 22468 38496 22520 38548
rect 3424 38360 3476 38412
rect 45192 38403 45244 38412
rect 45192 38369 45201 38403
rect 45201 38369 45235 38403
rect 45235 38369 45244 38403
rect 45192 38360 45244 38369
rect 21364 38335 21416 38344
rect 21364 38301 21373 38335
rect 21373 38301 21407 38335
rect 21407 38301 21416 38335
rect 21364 38292 21416 38301
rect 22008 38335 22060 38344
rect 22008 38301 22017 38335
rect 22017 38301 22051 38335
rect 22051 38301 22060 38335
rect 22008 38292 22060 38301
rect 23848 38335 23900 38344
rect 23848 38301 23857 38335
rect 23857 38301 23891 38335
rect 23891 38301 23900 38335
rect 23848 38292 23900 38301
rect 32312 38335 32364 38344
rect 32312 38301 32321 38335
rect 32321 38301 32355 38335
rect 32355 38301 32364 38335
rect 32312 38292 32364 38301
rect 51540 38335 51592 38344
rect 51540 38301 51549 38335
rect 51549 38301 51583 38335
rect 51583 38301 51592 38335
rect 51540 38292 51592 38301
rect 22652 38224 22704 38276
rect 33508 38224 33560 38276
rect 46848 38267 46900 38276
rect 46848 38233 46857 38267
rect 46857 38233 46891 38267
rect 46891 38233 46900 38267
rect 46848 38224 46900 38233
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 22652 37995 22704 38004
rect 22652 37961 22661 37995
rect 22661 37961 22695 37995
rect 22695 37961 22704 37995
rect 22652 37952 22704 37961
rect 33508 37995 33560 38004
rect 33508 37961 33517 37995
rect 33517 37961 33551 37995
rect 33551 37961 33560 37995
rect 33508 37952 33560 37961
rect 7196 37884 7248 37936
rect 28724 37884 28776 37936
rect 20628 37816 20680 37868
rect 22560 37859 22612 37868
rect 22560 37825 22569 37859
rect 22569 37825 22603 37859
rect 22603 37825 22612 37859
rect 22560 37816 22612 37825
rect 32312 37816 32364 37868
rect 28816 37748 28868 37800
rect 46388 37816 46440 37868
rect 48780 37859 48832 37868
rect 48780 37825 48789 37859
rect 48789 37825 48823 37859
rect 48823 37825 48832 37859
rect 48780 37816 48832 37825
rect 51172 37859 51224 37868
rect 51172 37825 51181 37859
rect 51181 37825 51215 37859
rect 51215 37825 51224 37859
rect 51172 37816 51224 37825
rect 48964 37748 49016 37800
rect 63408 37748 63460 37800
rect 6552 37612 6604 37664
rect 51264 37655 51316 37664
rect 51264 37621 51273 37655
rect 51273 37621 51307 37655
rect 51307 37621 51316 37655
rect 51264 37612 51316 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 4988 37272 5040 37324
rect 21364 37272 21416 37324
rect 51540 37272 51592 37324
rect 5264 37204 5316 37256
rect 6368 37204 6420 37256
rect 20628 37247 20680 37256
rect 20628 37213 20637 37247
rect 20637 37213 20671 37247
rect 20671 37213 20680 37247
rect 20628 37204 20680 37213
rect 22192 37204 22244 37256
rect 53380 37204 53432 37256
rect 20904 37179 20956 37188
rect 20904 37145 20913 37179
rect 20913 37145 20947 37179
rect 20947 37145 20956 37179
rect 20904 37136 20956 37145
rect 35440 37136 35492 37188
rect 51264 37136 51316 37188
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 6552 36839 6604 36848
rect 6552 36805 6561 36839
rect 6561 36805 6595 36839
rect 6595 36805 6604 36839
rect 6552 36796 6604 36805
rect 4988 36728 5040 36780
rect 6368 36771 6420 36780
rect 6368 36737 6377 36771
rect 6377 36737 6411 36771
rect 6411 36737 6420 36771
rect 6368 36728 6420 36737
rect 20628 36771 20680 36780
rect 20628 36737 20637 36771
rect 20637 36737 20671 36771
rect 20671 36737 20680 36771
rect 20628 36728 20680 36737
rect 38844 36771 38896 36780
rect 38844 36737 38853 36771
rect 38853 36737 38887 36771
rect 38887 36737 38896 36771
rect 38844 36728 38896 36737
rect 43904 36728 43956 36780
rect 4620 36660 4672 36712
rect 9772 36660 9824 36712
rect 34704 36660 34756 36712
rect 5448 36524 5500 36576
rect 38108 36524 38160 36576
rect 38936 36567 38988 36576
rect 38936 36533 38945 36567
rect 38945 36533 38979 36567
rect 38979 36533 38988 36567
rect 38936 36524 38988 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 20628 36320 20680 36372
rect 2872 36252 2924 36304
rect 5264 36227 5316 36236
rect 5264 36193 5273 36227
rect 5273 36193 5307 36227
rect 5307 36193 5316 36227
rect 5264 36184 5316 36193
rect 5448 36227 5500 36236
rect 5448 36193 5457 36227
rect 5457 36193 5491 36227
rect 5491 36193 5500 36227
rect 5448 36184 5500 36193
rect 31392 36116 31444 36168
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 38844 35776 38896 35828
rect 38936 35708 38988 35760
rect 38108 35683 38160 35692
rect 38108 35649 38117 35683
rect 38117 35649 38151 35683
rect 38151 35649 38160 35683
rect 38108 35640 38160 35649
rect 39764 35615 39816 35624
rect 39764 35581 39773 35615
rect 39773 35581 39807 35615
rect 39807 35581 39816 35615
rect 39764 35572 39816 35581
rect 63040 35615 63092 35624
rect 63040 35581 63049 35615
rect 63049 35581 63083 35615
rect 63083 35581 63092 35615
rect 63040 35572 63092 35581
rect 63776 35572 63828 35624
rect 66076 35572 66128 35624
rect 2780 35436 2832 35488
rect 4620 35436 4672 35488
rect 37096 35436 37148 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 63040 35232 63092 35284
rect 63776 35275 63828 35284
rect 63776 35241 63785 35275
rect 63785 35241 63819 35275
rect 63819 35241 63828 35275
rect 63776 35232 63828 35241
rect 3424 34892 3476 34944
rect 37096 35139 37148 35148
rect 37096 35105 37105 35139
rect 37105 35105 37139 35139
rect 37139 35105 37148 35139
rect 37096 35096 37148 35105
rect 63684 35071 63736 35080
rect 63684 35037 63693 35071
rect 63693 35037 63727 35071
rect 63727 35037 63736 35071
rect 63684 35028 63736 35037
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 42340 33940 42392 33992
rect 42892 33940 42944 33992
rect 42708 33915 42760 33924
rect 42708 33881 42717 33915
rect 42717 33881 42751 33915
rect 42751 33881 42760 33915
rect 42708 33872 42760 33881
rect 49056 33872 49108 33924
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 42340 33464 42392 33516
rect 42892 33507 42944 33516
rect 42892 33473 42901 33507
rect 42901 33473 42935 33507
rect 42935 33473 42944 33507
rect 42892 33464 42944 33473
rect 67456 33507 67508 33516
rect 67456 33473 67465 33507
rect 67465 33473 67499 33507
rect 67499 33473 67508 33507
rect 67456 33464 67508 33473
rect 41604 33439 41656 33448
rect 41604 33405 41613 33439
rect 41613 33405 41647 33439
rect 41647 33405 41656 33439
rect 41604 33396 41656 33405
rect 43076 33439 43128 33448
rect 43076 33405 43085 33439
rect 43085 33405 43119 33439
rect 43119 33405 43128 33439
rect 43076 33396 43128 33405
rect 65524 33396 65576 33448
rect 44088 33328 44140 33380
rect 62396 33303 62448 33312
rect 62396 33269 62405 33303
rect 62405 33269 62439 33303
rect 62439 33269 62448 33303
rect 62396 33260 62448 33269
rect 66444 33260 66496 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 43076 33056 43128 33108
rect 43812 32920 43864 32972
rect 42340 32852 42392 32904
rect 42984 32852 43036 32904
rect 44088 32895 44140 32904
rect 44088 32861 44097 32895
rect 44097 32861 44131 32895
rect 44131 32861 44140 32895
rect 51080 33056 51132 33108
rect 54208 33056 54260 33108
rect 62396 32920 62448 32972
rect 65800 32920 65852 32972
rect 44088 32852 44140 32861
rect 67456 32852 67508 32904
rect 61936 32784 61988 32836
rect 66168 32784 66220 32836
rect 44088 32716 44140 32768
rect 65984 32716 66036 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 61936 32555 61988 32564
rect 61936 32521 61945 32555
rect 61945 32521 61979 32555
rect 61979 32521 61988 32555
rect 61936 32512 61988 32521
rect 37372 32444 37424 32496
rect 44088 32487 44140 32496
rect 42340 32376 42392 32428
rect 44088 32453 44097 32487
rect 44097 32453 44131 32487
rect 44131 32453 44140 32487
rect 44088 32444 44140 32453
rect 65984 32487 66036 32496
rect 65984 32453 65993 32487
rect 65993 32453 66027 32487
rect 66027 32453 66036 32487
rect 65984 32444 66036 32453
rect 43812 32376 43864 32428
rect 60740 32376 60792 32428
rect 61844 32419 61896 32428
rect 61844 32385 61853 32419
rect 61853 32385 61887 32419
rect 61887 32385 61896 32419
rect 61844 32376 61896 32385
rect 65800 32419 65852 32428
rect 65800 32385 65809 32419
rect 65809 32385 65843 32419
rect 65843 32385 65852 32419
rect 65800 32376 65852 32385
rect 45468 32351 45520 32360
rect 45468 32317 45477 32351
rect 45477 32317 45511 32351
rect 45511 32317 45520 32351
rect 45468 32308 45520 32317
rect 67548 32351 67600 32360
rect 67548 32317 67557 32351
rect 67557 32317 67591 32351
rect 67591 32317 67600 32351
rect 67548 32308 67600 32317
rect 47584 32240 47636 32292
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 67640 31832 67692 31884
rect 67824 31875 67876 31884
rect 67824 31841 67833 31875
rect 67833 31841 67867 31875
rect 67867 31841 67876 31875
rect 67824 31832 67876 31841
rect 42708 31764 42760 31816
rect 66444 31739 66496 31748
rect 66444 31705 66453 31739
rect 66453 31705 66487 31739
rect 66487 31705 66496 31739
rect 66444 31696 66496 31705
rect 42616 31628 42668 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 42616 31399 42668 31408
rect 42616 31365 42625 31399
rect 42625 31365 42659 31399
rect 42659 31365 42668 31399
rect 42616 31356 42668 31365
rect 49056 31288 49108 31340
rect 67640 31331 67692 31340
rect 67640 31297 67649 31331
rect 67649 31297 67683 31331
rect 67683 31297 67692 31331
rect 67640 31288 67692 31297
rect 204 31220 256 31272
rect 59820 31220 59872 31272
rect 63132 31220 63184 31272
rect 42800 31084 42852 31136
rect 43352 31084 43404 31136
rect 51172 31084 51224 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 59820 30923 59872 30932
rect 59820 30889 59829 30923
rect 59829 30889 59863 30923
rect 59863 30889 59872 30923
rect 59820 30880 59872 30889
rect 22560 30744 22612 30796
rect 20628 30676 20680 30728
rect 26424 30719 26476 30728
rect 26424 30685 26433 30719
rect 26433 30685 26467 30719
rect 26467 30685 26476 30719
rect 26424 30676 26476 30685
rect 27068 30719 27120 30728
rect 27068 30685 27077 30719
rect 27077 30685 27111 30719
rect 27111 30685 27120 30719
rect 27068 30676 27120 30685
rect 28908 30651 28960 30660
rect 28908 30617 28917 30651
rect 28917 30617 28951 30651
rect 28951 30617 28960 30651
rect 28908 30608 28960 30617
rect 42340 30719 42392 30728
rect 42340 30685 42349 30719
rect 42349 30685 42383 30719
rect 42383 30685 42392 30719
rect 42340 30676 42392 30685
rect 42800 30608 42852 30660
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 42340 30268 42392 30320
rect 27068 30200 27120 30252
rect 8024 30175 8076 30184
rect 8024 30141 8033 30175
rect 8033 30141 8067 30175
rect 8067 30141 8076 30175
rect 8024 30132 8076 30141
rect 9036 30132 9088 30184
rect 4068 30064 4120 30116
rect 63132 30132 63184 30184
rect 66168 30132 66220 30184
rect 42984 30039 43036 30048
rect 42984 30005 42993 30039
rect 42993 30005 43027 30039
rect 43027 30005 43036 30039
rect 42984 29996 43036 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 8024 29792 8076 29844
rect 9036 29835 9088 29844
rect 9036 29801 9045 29835
rect 9045 29801 9079 29835
rect 9079 29801 9088 29835
rect 9036 29792 9088 29801
rect 3424 29656 3476 29708
rect 5632 29631 5684 29640
rect 5632 29597 5641 29631
rect 5641 29597 5675 29631
rect 5675 29597 5684 29631
rect 5632 29588 5684 29597
rect 9772 29588 9824 29640
rect 10784 29588 10836 29640
rect 12164 29588 12216 29640
rect 5448 29452 5500 29504
rect 20904 29656 20956 29708
rect 43628 29588 43680 29640
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 5632 29112 5684 29164
rect 12164 29155 12216 29164
rect 12164 29121 12173 29155
rect 12173 29121 12207 29155
rect 12207 29121 12216 29155
rect 12164 29112 12216 29121
rect 43628 29155 43680 29164
rect 43628 29121 43637 29155
rect 43637 29121 43671 29155
rect 43671 29121 43680 29155
rect 43628 29112 43680 29121
rect 12716 29044 12768 29096
rect 12808 29087 12860 29096
rect 12808 29053 12817 29087
rect 12817 29053 12851 29087
rect 12851 29053 12860 29087
rect 43812 29087 43864 29096
rect 12808 29044 12860 29053
rect 43812 29053 43821 29087
rect 43821 29053 43855 29087
rect 43855 29053 43864 29087
rect 43812 29044 43864 29053
rect 45192 29087 45244 29096
rect 45192 29053 45201 29087
rect 45201 29053 45235 29087
rect 45235 29053 45244 29087
rect 45192 29044 45244 29053
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 12716 28747 12768 28756
rect 12716 28713 12725 28747
rect 12725 28713 12759 28747
rect 12759 28713 12768 28747
rect 12716 28704 12768 28713
rect 43812 28704 43864 28756
rect 4988 28543 5040 28552
rect 4988 28509 4997 28543
rect 4997 28509 5031 28543
rect 5031 28509 5040 28543
rect 4988 28500 5040 28509
rect 5448 28543 5500 28552
rect 5448 28509 5457 28543
rect 5457 28509 5491 28543
rect 5491 28509 5500 28543
rect 5448 28500 5500 28509
rect 12624 28543 12676 28552
rect 12624 28509 12633 28543
rect 12633 28509 12667 28543
rect 12667 28509 12676 28543
rect 12624 28500 12676 28509
rect 43536 28543 43588 28552
rect 43536 28509 43545 28543
rect 43545 28509 43579 28543
rect 43579 28509 43588 28543
rect 43536 28500 43588 28509
rect 54208 28543 54260 28552
rect 54208 28509 54217 28543
rect 54217 28509 54251 28543
rect 54251 28509 54260 28543
rect 54208 28500 54260 28509
rect 54760 28500 54812 28552
rect 65524 28432 65576 28484
rect 5540 28407 5592 28416
rect 5540 28373 5549 28407
rect 5549 28373 5583 28407
rect 5583 28373 5592 28407
rect 5540 28364 5592 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 20628 28024 20680 28076
rect 41604 28024 41656 28076
rect 54760 28067 54812 28076
rect 54760 28033 54769 28067
rect 54769 28033 54803 28067
rect 54803 28033 54812 28067
rect 54760 28024 54812 28033
rect 9404 27820 9456 27872
rect 10324 27863 10376 27872
rect 10324 27829 10333 27863
rect 10333 27829 10367 27863
rect 10367 27829 10376 27863
rect 10324 27820 10376 27829
rect 26240 27863 26292 27872
rect 26240 27829 26249 27863
rect 26249 27829 26283 27863
rect 26283 27829 26292 27863
rect 27068 27863 27120 27872
rect 26240 27820 26292 27829
rect 27068 27829 27077 27863
rect 27077 27829 27111 27863
rect 27111 27829 27120 27863
rect 27068 27820 27120 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 3976 27548 4028 27600
rect 4988 27480 5040 27532
rect 5540 27480 5592 27532
rect 10324 27548 10376 27600
rect 23572 27548 23624 27600
rect 9404 27523 9456 27532
rect 9404 27489 9413 27523
rect 9413 27489 9447 27523
rect 9447 27489 9456 27523
rect 9404 27480 9456 27489
rect 9496 27480 9548 27532
rect 26240 27480 26292 27532
rect 4068 27276 4120 27328
rect 12808 27344 12860 27396
rect 27068 27344 27120 27396
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 8944 26256 8996 26308
rect 9496 26256 9548 26308
rect 4068 26188 4120 26240
rect 23572 26188 23624 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 34704 25891 34756 25900
rect 34704 25857 34713 25891
rect 34713 25857 34747 25891
rect 34747 25857 34756 25891
rect 34704 25848 34756 25857
rect 34796 25687 34848 25696
rect 34796 25653 34805 25687
rect 34805 25653 34839 25687
rect 34839 25653 34848 25687
rect 34796 25644 34848 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 34796 25304 34848 25356
rect 34888 25279 34940 25288
rect 34888 25245 34897 25279
rect 34897 25245 34931 25279
rect 34931 25245 34940 25279
rect 34888 25236 34940 25245
rect 36728 25211 36780 25220
rect 36728 25177 36737 25211
rect 36737 25177 36771 25211
rect 36771 25177 36780 25211
rect 36728 25168 36780 25177
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 28816 24803 28868 24812
rect 28816 24769 28825 24803
rect 28825 24769 28859 24803
rect 28859 24769 28868 24803
rect 28816 24760 28868 24769
rect 34888 24760 34940 24812
rect 28356 24599 28408 24608
rect 28356 24565 28365 24599
rect 28365 24565 28399 24599
rect 28399 24565 28408 24599
rect 28356 24556 28408 24565
rect 28540 24556 28592 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 58164 24148 58216 24200
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 28540 23783 28592 23792
rect 28540 23749 28549 23783
rect 28549 23749 28583 23783
rect 28583 23749 28592 23783
rect 28540 23740 28592 23749
rect 28356 23715 28408 23724
rect 28356 23681 28365 23715
rect 28365 23681 28399 23715
rect 28399 23681 28408 23715
rect 28356 23672 28408 23681
rect 58164 23715 58216 23724
rect 58164 23681 58173 23715
rect 58173 23681 58207 23715
rect 58207 23681 58216 23715
rect 58164 23672 58216 23681
rect 6920 23604 6972 23656
rect 58348 23647 58400 23656
rect 58348 23613 58357 23647
rect 58357 23613 58391 23647
rect 58391 23613 58400 23647
rect 58348 23604 58400 23613
rect 65984 23604 66036 23656
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 36728 23264 36780 23316
rect 58348 23264 58400 23316
rect 66168 23196 66220 23248
rect 10784 23103 10836 23112
rect 10784 23069 10793 23103
rect 10793 23069 10827 23103
rect 10827 23069 10836 23103
rect 10784 23060 10836 23069
rect 11612 23103 11664 23112
rect 11612 23069 11621 23103
rect 11621 23069 11655 23103
rect 11655 23069 11664 23103
rect 11612 23060 11664 23069
rect 57888 23103 57940 23112
rect 57888 23069 57897 23103
rect 57897 23069 57931 23103
rect 57931 23069 57940 23103
rect 57888 23060 57940 23069
rect 60740 23103 60792 23112
rect 60740 23069 60749 23103
rect 60749 23069 60783 23103
rect 60783 23069 60792 23103
rect 60740 23060 60792 23069
rect 60648 22992 60700 23044
rect 10784 22924 10836 22976
rect 60832 22967 60884 22976
rect 60832 22933 60841 22967
rect 60841 22933 60875 22967
rect 60875 22933 60884 22967
rect 60832 22924 60884 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 60832 22695 60884 22704
rect 60832 22661 60841 22695
rect 60841 22661 60875 22695
rect 60875 22661 60884 22695
rect 60832 22652 60884 22661
rect 47584 22584 47636 22636
rect 57888 22584 57940 22636
rect 60648 22627 60700 22636
rect 60648 22593 60657 22627
rect 60657 22593 60691 22627
rect 60691 22593 60700 22627
rect 60648 22584 60700 22593
rect 62488 22559 62540 22568
rect 62488 22525 62497 22559
rect 62497 22525 62531 22559
rect 62531 22525 62540 22559
rect 62488 22516 62540 22525
rect 4712 22423 4764 22432
rect 4712 22389 4721 22423
rect 4721 22389 4755 22423
rect 4755 22389 4764 22423
rect 4712 22380 4764 22389
rect 50528 22380 50580 22432
rect 51356 22423 51408 22432
rect 51356 22389 51365 22423
rect 51365 22389 51399 22423
rect 51399 22389 51408 22423
rect 51356 22380 51408 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 3332 22108 3384 22160
rect 4712 22040 4764 22092
rect 10784 22083 10836 22092
rect 10784 22049 10793 22083
rect 10793 22049 10827 22083
rect 10827 22049 10836 22083
rect 10784 22040 10836 22049
rect 12348 22083 12400 22092
rect 12348 22049 12357 22083
rect 12357 22049 12391 22083
rect 12391 22049 12400 22083
rect 12348 22040 12400 22049
rect 50528 22083 50580 22092
rect 50528 22049 50537 22083
rect 50537 22049 50571 22083
rect 50571 22049 50580 22083
rect 50528 22040 50580 22049
rect 50804 22083 50856 22092
rect 50804 22049 50813 22083
rect 50813 22049 50847 22083
rect 50847 22049 50856 22083
rect 50804 22040 50856 22049
rect 62948 22015 63000 22024
rect 5080 21904 5132 21956
rect 11612 21904 11664 21956
rect 62948 21981 62957 22015
rect 62957 21981 62991 22015
rect 62991 21981 63000 22015
rect 62948 21972 63000 21981
rect 51356 21904 51408 21956
rect 63316 21836 63368 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 5080 21675 5132 21684
rect 5080 21641 5089 21675
rect 5089 21641 5123 21675
rect 5123 21641 5132 21675
rect 5080 21632 5132 21641
rect 63316 21607 63368 21616
rect 63316 21573 63325 21607
rect 63325 21573 63359 21607
rect 63359 21573 63368 21607
rect 63316 21564 63368 21573
rect 4896 21496 4948 21548
rect 63132 21471 63184 21480
rect 63132 21437 63141 21471
rect 63141 21437 63175 21471
rect 63175 21437 63184 21471
rect 63132 21428 63184 21437
rect 66076 21428 66128 21480
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 63132 21088 63184 21140
rect 49792 20748 49844 20800
rect 50804 20748 50856 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 32128 19796 32180 19848
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 3516 19388 3568 19440
rect 32128 19363 32180 19372
rect 32128 19329 32137 19363
rect 32137 19329 32171 19363
rect 32171 19329 32180 19363
rect 32128 19320 32180 19329
rect 32312 19295 32364 19304
rect 32312 19261 32321 19295
rect 32321 19261 32355 19295
rect 32355 19261 32364 19295
rect 32312 19252 32364 19261
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 32312 18912 32364 18964
rect 45376 18708 45428 18760
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 5448 18071 5500 18080
rect 5448 18037 5457 18071
rect 5457 18037 5491 18071
rect 5491 18037 5500 18071
rect 5448 18028 5500 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 5448 17688 5500 17740
rect 6828 17731 6880 17740
rect 6828 17697 6837 17731
rect 6837 17697 6871 17731
rect 6871 17697 6880 17731
rect 6828 17688 6880 17697
rect 62948 17620 63000 17672
rect 63040 17620 63092 17672
rect 5540 17552 5592 17604
rect 63224 17484 63276 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 5540 17323 5592 17332
rect 5540 17289 5549 17323
rect 5549 17289 5583 17323
rect 5583 17289 5592 17323
rect 5540 17280 5592 17289
rect 63224 17255 63276 17264
rect 63224 17221 63233 17255
rect 63233 17221 63267 17255
rect 63267 17221 63276 17255
rect 63224 17212 63276 17221
rect 4896 17144 4948 17196
rect 5448 17187 5500 17196
rect 5448 17153 5457 17187
rect 5457 17153 5491 17187
rect 5491 17153 5500 17187
rect 5448 17144 5500 17153
rect 63040 17187 63092 17196
rect 63040 17153 63049 17187
rect 63049 17153 63083 17187
rect 63083 17153 63092 17187
rect 63040 17144 63092 17153
rect 64788 17119 64840 17128
rect 64788 17085 64797 17119
rect 64797 17085 64831 17119
rect 64831 17085 64840 17119
rect 64788 17076 64840 17085
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 3332 16532 3384 16584
rect 8944 16532 8996 16584
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 12808 15444 12860 15496
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 62488 15104 62540 15156
rect 66076 15104 66128 15156
rect 12808 15011 12860 15020
rect 12808 14977 12817 15011
rect 12817 14977 12851 15011
rect 12851 14977 12860 15011
rect 12808 14968 12860 14977
rect 12992 14943 13044 14952
rect 12992 14909 13001 14943
rect 13001 14909 13035 14943
rect 13035 14909 13044 14943
rect 12992 14900 13044 14909
rect 13544 14943 13596 14952
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 12992 14560 13044 14612
rect 5448 14356 5500 14408
rect 19432 14356 19484 14408
rect 22100 14399 22152 14408
rect 22100 14365 22109 14399
rect 22109 14365 22143 14399
rect 22143 14365 22152 14399
rect 22100 14356 22152 14365
rect 22192 14263 22244 14272
rect 22192 14229 22201 14263
rect 22201 14229 22235 14263
rect 22235 14229 22244 14263
rect 22192 14220 22244 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 22192 13991 22244 14000
rect 22192 13957 22201 13991
rect 22201 13957 22235 13991
rect 22235 13957 22244 13991
rect 22192 13948 22244 13957
rect 19432 13923 19484 13932
rect 19432 13889 19441 13923
rect 19441 13889 19475 13923
rect 19475 13889 19484 13923
rect 19432 13880 19484 13889
rect 19616 13855 19668 13864
rect 19616 13821 19625 13855
rect 19625 13821 19659 13855
rect 19659 13821 19668 13855
rect 19616 13812 19668 13821
rect 3332 13744 3384 13796
rect 22192 13812 22244 13864
rect 22560 13855 22612 13864
rect 22560 13821 22569 13855
rect 22569 13821 22603 13855
rect 22603 13821 22612 13855
rect 22560 13812 22612 13821
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 19616 13472 19668 13524
rect 22192 13515 22244 13524
rect 22192 13481 22201 13515
rect 22201 13481 22235 13515
rect 22235 13481 22244 13515
rect 22192 13472 22244 13481
rect 22100 13268 22152 13320
rect 35624 13175 35676 13184
rect 35624 13141 35633 13175
rect 35633 13141 35667 13175
rect 35667 13141 35676 13175
rect 35624 13132 35676 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 35440 12588 35492 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 26884 12180 26936 12232
rect 45284 12316 45336 12368
rect 35440 12291 35492 12300
rect 35440 12257 35449 12291
rect 35449 12257 35483 12291
rect 35483 12257 35492 12291
rect 35440 12248 35492 12257
rect 35624 12291 35676 12300
rect 35624 12257 35633 12291
rect 35633 12257 35667 12291
rect 35667 12257 35676 12291
rect 35624 12248 35676 12257
rect 36084 12291 36136 12300
rect 36084 12257 36093 12291
rect 36093 12257 36127 12291
rect 36127 12257 36136 12291
rect 36084 12248 36136 12257
rect 63408 12180 63460 12232
rect 34428 12044 34480 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 34428 11815 34480 11824
rect 34428 11781 34437 11815
rect 34437 11781 34471 11815
rect 34471 11781 34480 11815
rect 34428 11772 34480 11781
rect 63408 11747 63460 11756
rect 63408 11713 63417 11747
rect 63417 11713 63451 11747
rect 63451 11713 63460 11747
rect 63408 11704 63460 11713
rect 34796 11679 34848 11688
rect 34796 11645 34805 11679
rect 34805 11645 34839 11679
rect 34839 11645 34848 11679
rect 34796 11636 34848 11645
rect 63316 11636 63368 11688
rect 65248 11679 65300 11688
rect 65248 11645 65257 11679
rect 65257 11645 65291 11679
rect 65291 11645 65300 11679
rect 65248 11636 65300 11645
rect 24584 11500 24636 11552
rect 30104 11500 30156 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 63316 11339 63368 11348
rect 63316 11305 63325 11339
rect 63325 11305 63359 11339
rect 63359 11305 63368 11339
rect 63316 11296 63368 11305
rect 5816 11228 5868 11280
rect 3608 11160 3660 11212
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 26884 11135 26936 11144
rect 26884 11101 26893 11135
rect 26893 11101 26927 11135
rect 26927 11101 26936 11135
rect 26884 11092 26936 11101
rect 30104 11135 30156 11144
rect 30104 11101 30113 11135
rect 30113 11101 30147 11135
rect 30147 11101 30156 11135
rect 30104 11092 30156 11101
rect 63684 11092 63736 11144
rect 19984 11024 20036 11076
rect 24768 11067 24820 11076
rect 24768 11033 24777 11067
rect 24777 11033 24811 11067
rect 24811 11033 24820 11067
rect 24768 11024 24820 11033
rect 30656 11024 30708 11076
rect 35072 11067 35124 11076
rect 35072 11033 35081 11067
rect 35081 11033 35115 11067
rect 35115 11033 35124 11067
rect 35072 11024 35124 11033
rect 26240 10956 26292 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 24860 10752 24912 10804
rect 30656 10795 30708 10804
rect 30656 10761 30665 10795
rect 30665 10761 30699 10795
rect 30699 10761 30708 10795
rect 30656 10752 30708 10761
rect 35072 10752 35124 10804
rect 26884 10616 26936 10668
rect 48964 10616 49016 10668
rect 26056 10412 26108 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 26056 10115 26108 10124
rect 26056 10081 26065 10115
rect 26065 10081 26099 10115
rect 26099 10081 26108 10115
rect 26056 10072 26108 10081
rect 26240 10115 26292 10124
rect 26240 10081 26249 10115
rect 26249 10081 26283 10115
rect 26283 10081 26292 10115
rect 26240 10072 26292 10081
rect 43352 10047 43404 10056
rect 43352 10013 43361 10047
rect 43361 10013 43395 10047
rect 43395 10013 43404 10047
rect 43352 10004 43404 10013
rect 54392 10004 54444 10056
rect 27804 9936 27856 9988
rect 43444 9911 43496 9920
rect 43444 9877 43453 9911
rect 43453 9877 43487 9911
rect 43487 9877 43496 9911
rect 43444 9868 43496 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 43444 9639 43496 9648
rect 43444 9605 43453 9639
rect 43453 9605 43487 9639
rect 43487 9605 43496 9639
rect 43444 9596 43496 9605
rect 43536 9460 43588 9512
rect 43812 9503 43864 9512
rect 43812 9469 43821 9503
rect 43821 9469 43855 9503
rect 43855 9469 43864 9503
rect 43812 9460 43864 9469
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 43536 9163 43588 9172
rect 43536 9129 43545 9163
rect 43545 9129 43579 9163
rect 43579 9129 43588 9163
rect 43536 9120 43588 9129
rect 20 8848 72 8900
rect 54392 8959 54444 8968
rect 54392 8925 54401 8959
rect 54401 8925 54435 8959
rect 54435 8925 54444 8959
rect 54392 8916 54444 8925
rect 54760 8916 54812 8968
rect 27068 8848 27120 8900
rect 54944 8780 54996 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 27068 8619 27120 8628
rect 27068 8585 27077 8619
rect 27077 8585 27111 8619
rect 27111 8585 27120 8619
rect 27068 8576 27120 8585
rect 54944 8551 54996 8560
rect 54944 8517 54953 8551
rect 54953 8517 54987 8551
rect 54987 8517 54996 8551
rect 54944 8508 54996 8517
rect 43352 8440 43404 8492
rect 54760 8483 54812 8492
rect 54760 8449 54769 8483
rect 54769 8449 54803 8483
rect 54803 8449 54812 8483
rect 54760 8440 54812 8449
rect 59268 8372 59320 8424
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 45192 4088 45244 4140
rect 47032 4088 47084 4140
rect 45100 4020 45152 4072
rect 46848 4020 46900 4072
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 24492 3544 24544 3596
rect 28908 3544 28960 3596
rect 68928 3544 68980 3596
rect 4620 3476 4672 3528
rect 6828 3476 6880 3528
rect 10968 3476 11020 3528
rect 12348 3476 12400 3528
rect 26424 3476 26476 3528
rect 40684 3519 40736 3528
rect 40684 3485 40693 3519
rect 40693 3485 40727 3519
rect 40727 3485 40736 3519
rect 40684 3476 40736 3485
rect 67824 3476 67876 3528
rect 69572 3476 69624 3528
rect 27068 3451 27120 3460
rect 27068 3417 27077 3451
rect 27077 3417 27111 3451
rect 27111 3417 27120 3451
rect 27068 3408 27120 3417
rect 41788 3408 41840 3460
rect 41236 3340 41288 3392
rect 45468 3408 45520 3460
rect 61200 3408 61252 3460
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 41788 3179 41840 3188
rect 41788 3145 41797 3179
rect 41797 3145 41831 3179
rect 41831 3145 41840 3179
rect 41788 3136 41840 3145
rect 56508 3136 56560 3188
rect 62488 3136 62540 3188
rect 26424 3043 26476 3052
rect 26424 3009 26433 3043
rect 26433 3009 26467 3043
rect 26467 3009 26476 3043
rect 26424 3000 26476 3009
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 41696 3043 41748 3052
rect 41696 3009 41705 3043
rect 41705 3009 41739 3043
rect 41739 3009 41748 3043
rect 41696 3000 41748 3009
rect 42984 3000 43036 3052
rect 27620 2975 27672 2984
rect 27620 2941 27629 2975
rect 27629 2941 27663 2975
rect 27663 2941 27672 2975
rect 27620 2932 27672 2941
rect 39580 2975 39632 2984
rect 14832 2864 14884 2916
rect 39580 2941 39589 2975
rect 39589 2941 39623 2975
rect 39623 2941 39632 2975
rect 39580 2932 39632 2941
rect 39948 2975 40000 2984
rect 39948 2941 39957 2975
rect 39957 2941 39991 2975
rect 39991 2941 40000 2975
rect 39948 2932 40000 2941
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 27068 2592 27120 2644
rect 27620 2592 27672 2644
rect 39580 2592 39632 2644
rect 40684 2592 40736 2644
rect 26976 2388 27028 2440
rect 41696 2388 41748 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 3424 1300 3476 1352
rect 27804 1300 27856 1352
rect 59268 1300 59320 1352
rect 66168 1300 66220 1352
<< metal2 >>
rect 634 71200 746 72000
rect 1278 71200 1390 72000
rect 1490 71496 1546 71505
rect 1490 71431 1546 71440
rect 1504 69426 1532 71431
rect 2566 71200 2678 72000
rect 3854 71200 3966 72000
rect 5142 71346 5254 72000
rect 4632 71318 5254 71346
rect 1492 69420 1544 69426
rect 1492 69362 1544 69368
rect 3514 68776 3570 68785
rect 3514 68711 3570 68720
rect 3422 67416 3478 67425
rect 3422 67351 3478 67360
rect 1400 60648 1452 60654
rect 1398 60616 1400 60625
rect 1452 60616 1454 60625
rect 1398 60551 1454 60560
rect 3330 59256 3386 59265
rect 3330 59191 3386 59200
rect 3344 58954 3372 59191
rect 3332 58948 3384 58954
rect 3332 58890 3384 58896
rect 2964 55616 3016 55622
rect 2964 55558 3016 55564
rect 2976 55214 3004 55558
rect 2884 55186 3004 55214
rect 2778 55176 2834 55185
rect 2778 55111 2834 55120
rect 2792 54058 2820 55111
rect 2780 54052 2832 54058
rect 2780 53994 2832 54000
rect 2884 51105 2912 55186
rect 3330 53816 3386 53825
rect 3330 53751 3386 53760
rect 2962 52456 3018 52465
rect 2962 52391 3018 52400
rect 2976 52086 3004 52391
rect 2964 52080 3016 52086
rect 2964 52022 3016 52028
rect 2870 51096 2926 51105
rect 2870 51031 2926 51040
rect 3344 50998 3372 53751
rect 3332 50992 3384 50998
rect 3332 50934 3384 50940
rect 3436 45014 3464 67351
rect 3528 53650 3556 68711
rect 3896 68134 3924 71200
rect 4214 69116 4522 69125
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69051 4522 69060
rect 3884 68128 3936 68134
rect 3884 68070 3936 68076
rect 4214 68028 4522 68037
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67963 4522 67972
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 4632 64530 4660 71318
rect 5142 71200 5254 71318
rect 6430 71200 6542 72000
rect 7718 71200 7830 72000
rect 9006 71200 9118 72000
rect 10294 71200 10406 72000
rect 11582 71346 11694 72000
rect 11072 71318 11694 71346
rect 6472 68406 6500 71200
rect 6460 68400 6512 68406
rect 6460 68342 6512 68348
rect 5540 68128 5592 68134
rect 5540 68070 5592 68076
rect 5552 64938 5580 68070
rect 6736 65544 6788 65550
rect 6736 65486 6788 65492
rect 6748 65074 6776 65486
rect 6736 65068 6788 65074
rect 6736 65010 6788 65016
rect 6920 65000 6972 65006
rect 6920 64942 6972 64948
rect 5540 64932 5592 64938
rect 5540 64874 5592 64880
rect 6932 64666 6960 64942
rect 6920 64660 6972 64666
rect 6920 64602 6972 64608
rect 4620 64524 4672 64530
rect 4620 64466 4672 64472
rect 7196 64456 7248 64462
rect 7196 64398 7248 64404
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 5724 54052 5776 54058
rect 5724 53994 5776 54000
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 3516 53644 3568 53650
rect 3516 53586 3568 53592
rect 5264 52896 5316 52902
rect 5264 52838 5316 52844
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 5276 52562 5304 52838
rect 5736 52562 5764 53994
rect 5264 52556 5316 52562
rect 5264 52498 5316 52504
rect 5632 52556 5684 52562
rect 5632 52498 5684 52504
rect 5724 52556 5776 52562
rect 5724 52498 5776 52504
rect 5644 52154 5672 52498
rect 5632 52148 5684 52154
rect 5632 52090 5684 52096
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 6920 50312 6972 50318
rect 6920 50254 6972 50260
rect 6932 49842 6960 50254
rect 6920 49836 6972 49842
rect 6920 49778 6972 49784
rect 4068 49768 4120 49774
rect 4066 49736 4068 49745
rect 7104 49768 7156 49774
rect 4120 49736 4122 49745
rect 7104 49710 7156 49716
rect 4066 49671 4122 49680
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 7116 49434 7144 49710
rect 7104 49428 7156 49434
rect 7104 49370 7156 49376
rect 7208 49230 7236 64398
rect 11072 56914 11100 71318
rect 11582 71200 11694 71318
rect 12870 71200 12982 72000
rect 14158 71200 14270 72000
rect 15446 71200 15558 72000
rect 16734 71200 16846 72000
rect 18022 71200 18134 72000
rect 19310 71200 19422 72000
rect 20598 71200 20710 72000
rect 21886 71200 21998 72000
rect 23174 71200 23286 72000
rect 23818 71200 23930 72000
rect 25106 71200 25218 72000
rect 26394 71200 26506 72000
rect 27682 71346 27794 72000
rect 28970 71346 29082 72000
rect 27682 71318 28856 71346
rect 27682 71200 27794 71318
rect 16776 68474 16804 71200
rect 19574 69660 19882 69669
rect 19574 69658 19580 69660
rect 19636 69658 19660 69660
rect 19716 69658 19740 69660
rect 19796 69658 19820 69660
rect 19876 69658 19882 69660
rect 19636 69606 19638 69658
rect 19818 69606 19820 69658
rect 19574 69604 19580 69606
rect 19636 69604 19660 69606
rect 19716 69604 19740 69606
rect 19796 69604 19820 69606
rect 19876 69604 19882 69606
rect 19574 69595 19882 69604
rect 19574 68572 19882 68581
rect 19574 68570 19580 68572
rect 19636 68570 19660 68572
rect 19716 68570 19740 68572
rect 19796 68570 19820 68572
rect 19876 68570 19882 68572
rect 19636 68518 19638 68570
rect 19818 68518 19820 68570
rect 19574 68516 19580 68518
rect 19636 68516 19660 68518
rect 19716 68516 19740 68518
rect 19796 68516 19820 68518
rect 19876 68516 19882 68518
rect 19574 68507 19882 68516
rect 16764 68468 16816 68474
rect 16764 68410 16816 68416
rect 22744 68400 22796 68406
rect 22744 68342 22796 68348
rect 19574 67484 19882 67493
rect 19574 67482 19580 67484
rect 19636 67482 19660 67484
rect 19716 67482 19740 67484
rect 19796 67482 19820 67484
rect 19876 67482 19882 67484
rect 19636 67430 19638 67482
rect 19818 67430 19820 67482
rect 19574 67428 19580 67430
rect 19636 67428 19660 67430
rect 19716 67428 19740 67430
rect 19796 67428 19820 67430
rect 19876 67428 19882 67430
rect 19574 67419 19882 67428
rect 19574 66396 19882 66405
rect 19574 66394 19580 66396
rect 19636 66394 19660 66396
rect 19716 66394 19740 66396
rect 19796 66394 19820 66396
rect 19876 66394 19882 66396
rect 19636 66342 19638 66394
rect 19818 66342 19820 66394
rect 19574 66340 19580 66342
rect 19636 66340 19660 66342
rect 19716 66340 19740 66342
rect 19796 66340 19820 66342
rect 19876 66340 19882 66342
rect 19574 66331 19882 66340
rect 19574 65308 19882 65317
rect 19574 65306 19580 65308
rect 19636 65306 19660 65308
rect 19716 65306 19740 65308
rect 19796 65306 19820 65308
rect 19876 65306 19882 65308
rect 19636 65254 19638 65306
rect 19818 65254 19820 65306
rect 19574 65252 19580 65254
rect 19636 65252 19660 65254
rect 19716 65252 19740 65254
rect 19796 65252 19820 65254
rect 19876 65252 19882 65254
rect 19574 65243 19882 65252
rect 19574 64220 19882 64229
rect 19574 64218 19580 64220
rect 19636 64218 19660 64220
rect 19716 64218 19740 64220
rect 19796 64218 19820 64220
rect 19876 64218 19882 64220
rect 19636 64166 19638 64218
rect 19818 64166 19820 64218
rect 19574 64164 19580 64166
rect 19636 64164 19660 64166
rect 19716 64164 19740 64166
rect 19796 64164 19820 64166
rect 19876 64164 19882 64166
rect 19574 64155 19882 64164
rect 19574 63132 19882 63141
rect 19574 63130 19580 63132
rect 19636 63130 19660 63132
rect 19716 63130 19740 63132
rect 19796 63130 19820 63132
rect 19876 63130 19882 63132
rect 19636 63078 19638 63130
rect 19818 63078 19820 63130
rect 19574 63076 19580 63078
rect 19636 63076 19660 63078
rect 19716 63076 19740 63078
rect 19796 63076 19820 63078
rect 19876 63076 19882 63078
rect 19574 63067 19882 63076
rect 19574 62044 19882 62053
rect 19574 62042 19580 62044
rect 19636 62042 19660 62044
rect 19716 62042 19740 62044
rect 19796 62042 19820 62044
rect 19876 62042 19882 62044
rect 19636 61990 19638 62042
rect 19818 61990 19820 62042
rect 19574 61988 19580 61990
rect 19636 61988 19660 61990
rect 19716 61988 19740 61990
rect 19796 61988 19820 61990
rect 19876 61988 19882 61990
rect 19574 61979 19882 61988
rect 19574 60956 19882 60965
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60891 19882 60900
rect 22756 60518 22784 68342
rect 23216 68338 23244 71200
rect 25148 69018 25176 71200
rect 25136 69012 25188 69018
rect 25136 68954 25188 68960
rect 28264 69012 28316 69018
rect 28264 68954 28316 68960
rect 24124 68400 24176 68406
rect 24124 68342 24176 68348
rect 23204 68332 23256 68338
rect 23204 68274 23256 68280
rect 23020 61192 23072 61198
rect 23020 61134 23072 61140
rect 23032 60722 23060 61134
rect 23020 60716 23072 60722
rect 23020 60658 23072 60664
rect 23400 60710 23704 60738
rect 23400 60518 23428 60710
rect 23676 60654 23704 60710
rect 23572 60648 23624 60654
rect 23572 60590 23624 60596
rect 23664 60648 23716 60654
rect 23664 60590 23716 60596
rect 22744 60512 22796 60518
rect 22744 60454 22796 60460
rect 23388 60512 23440 60518
rect 23388 60454 23440 60460
rect 23584 60314 23612 60590
rect 23572 60308 23624 60314
rect 23572 60250 23624 60256
rect 19574 59868 19882 59877
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59803 19882 59812
rect 19574 58780 19882 58789
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58715 19882 58724
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 11060 56908 11112 56914
rect 11060 56850 11112 56856
rect 11336 56772 11388 56778
rect 11336 56714 11388 56720
rect 11348 56506 11376 56714
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 11336 56500 11388 56506
rect 11336 56442 11388 56448
rect 20628 56500 20680 56506
rect 20628 56442 20680 56448
rect 20640 56370 20668 56442
rect 11520 56364 11572 56370
rect 11520 56306 11572 56312
rect 20628 56364 20680 56370
rect 20628 56306 20680 56312
rect 7564 52896 7616 52902
rect 7564 52838 7616 52844
rect 7576 52018 7604 52838
rect 11532 52494 11560 56306
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 11520 52488 11572 52494
rect 11520 52430 11572 52436
rect 7748 52352 7800 52358
rect 7748 52294 7800 52300
rect 7760 52086 7788 52294
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 7748 52080 7800 52086
rect 7748 52022 7800 52028
rect 7564 52012 7616 52018
rect 7564 51954 7616 51960
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 7196 49224 7248 49230
rect 7196 49166 7248 49172
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4066 47696 4122 47705
rect 4066 47631 4122 47640
rect 4080 47598 4108 47631
rect 4068 47592 4120 47598
rect 4068 47534 4120 47540
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 3424 45008 3476 45014
rect 3424 44950 3476 44956
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 3054 40896 3110 40905
rect 3054 40831 3110 40840
rect 3068 40118 3096 40831
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 3056 40112 3108 40118
rect 3056 40054 3108 40060
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 3330 39536 3386 39545
rect 3330 39471 3386 39480
rect 3344 39370 3372 39471
rect 3332 39364 3384 39370
rect 3332 39306 3384 39312
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 3424 38412 3476 38418
rect 3424 38354 3476 38360
rect 3436 38185 3464 38354
rect 3422 38176 3478 38185
rect 3422 38111 3478 38120
rect 7208 37942 7236 49166
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 14740 45280 14792 45286
rect 14740 45222 14792 45228
rect 14752 44946 14780 45222
rect 14740 44940 14792 44946
rect 14740 44882 14792 44888
rect 15108 44804 15160 44810
rect 15108 44746 15160 44752
rect 15120 44538 15148 44746
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 15108 44532 15160 44538
rect 15108 44474 15160 44480
rect 13728 44396 13780 44402
rect 13728 44338 13780 44344
rect 13740 42226 13768 44338
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 12624 42220 12676 42226
rect 12624 42162 12676 42168
rect 13728 42220 13780 42226
rect 13728 42162 13780 42168
rect 9588 39840 9640 39846
rect 9588 39782 9640 39788
rect 9600 39506 9628 39782
rect 9588 39500 9640 39506
rect 9588 39442 9640 39448
rect 9864 39364 9916 39370
rect 9864 39306 9916 39312
rect 9876 39098 9904 39306
rect 9864 39092 9916 39098
rect 9864 39034 9916 39040
rect 9772 38956 9824 38962
rect 9772 38898 9824 38904
rect 7196 37936 7248 37942
rect 7196 37878 7248 37884
rect 6552 37664 6604 37670
rect 6552 37606 6604 37612
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4988 37324 5040 37330
rect 4988 37266 5040 37272
rect 2870 36816 2926 36825
rect 5000 36786 5028 37266
rect 5264 37256 5316 37262
rect 5264 37198 5316 37204
rect 6368 37256 6420 37262
rect 6368 37198 6420 37204
rect 2870 36751 2926 36760
rect 4988 36780 5040 36786
rect 2884 36310 2912 36751
rect 4988 36722 5040 36728
rect 4620 36712 4672 36718
rect 4620 36654 4672 36660
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 2872 36304 2924 36310
rect 2872 36246 2924 36252
rect 4632 35494 4660 36654
rect 5000 35894 5028 36722
rect 5276 36242 5304 37198
rect 6380 36786 6408 37198
rect 6564 36854 6592 37606
rect 6552 36848 6604 36854
rect 6552 36790 6604 36796
rect 6368 36780 6420 36786
rect 6368 36722 6420 36728
rect 9784 36718 9812 38898
rect 9772 36712 9824 36718
rect 9772 36654 9824 36660
rect 5448 36576 5500 36582
rect 5448 36518 5500 36524
rect 5460 36242 5488 36518
rect 5264 36236 5316 36242
rect 5264 36178 5316 36184
rect 5448 36236 5500 36242
rect 5448 36178 5500 36184
rect 4908 35866 5028 35894
rect 2780 35488 2832 35494
rect 2778 35456 2780 35465
rect 4620 35488 4672 35494
rect 2832 35456 2834 35465
rect 4620 35430 4672 35436
rect 2778 35391 2834 35400
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 3424 34944 3476 34950
rect 3424 34886 3476 34892
rect 3436 31385 3464 34886
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3422 31376 3478 31385
rect 3422 31311 3478 31320
rect 204 31272 256 31278
rect 204 31214 256 31220
rect 216 16574 244 31214
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4068 30116 4120 30122
rect 4068 30058 4120 30064
rect 4080 30025 4108 30058
rect 4066 30016 4122 30025
rect 4066 29951 4122 29960
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3424 29708 3476 29714
rect 3424 29650 3476 29656
rect 3330 22536 3386 22545
rect 3330 22471 3386 22480
rect 3344 22166 3372 22471
rect 3332 22160 3384 22166
rect 3332 22102 3384 22108
rect 3332 16584 3384 16590
rect 216 16546 704 16574
rect 20 8900 72 8906
rect 20 8842 72 8848
rect 32 800 60 8842
rect 676 800 704 16546
rect 3332 16526 3384 16532
rect 3344 15745 3372 16526
rect 3330 15736 3386 15745
rect 3330 15671 3386 15680
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 3344 13025 3372 13738
rect 3330 13016 3386 13025
rect 3330 12951 3386 12960
rect 3436 3505 3464 29650
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3976 27600 4028 27606
rect 3976 27542 4028 27548
rect 3988 23905 4016 27542
rect 4068 27328 4120 27334
rect 4066 27296 4068 27305
rect 4120 27296 4122 27305
rect 4066 27231 4122 27240
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4068 26240 4120 26246
rect 4068 26182 4120 26188
rect 4080 25945 4108 26182
rect 4066 25936 4122 25945
rect 4066 25871 4122 25880
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3974 23896 4030 23905
rect 3974 23831 4030 23840
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4724 22098 4752 22374
rect 4712 22092 4764 22098
rect 4712 22034 4764 22040
rect 4908 21554 4936 35866
rect 8024 30184 8076 30190
rect 8024 30126 8076 30132
rect 9036 30184 9088 30190
rect 9036 30126 9088 30132
rect 8036 29850 8064 30126
rect 9048 29850 9076 30126
rect 8024 29844 8076 29850
rect 8024 29786 8076 29792
rect 9036 29844 9088 29850
rect 9036 29786 9088 29792
rect 9784 29646 9812 36654
rect 5632 29640 5684 29646
rect 5632 29582 5684 29588
rect 9772 29640 9824 29646
rect 9772 29582 9824 29588
rect 10784 29640 10836 29646
rect 10784 29582 10836 29588
rect 12164 29640 12216 29646
rect 12164 29582 12216 29588
rect 5448 29504 5500 29510
rect 5448 29446 5500 29452
rect 5460 28558 5488 29446
rect 5644 29170 5672 29582
rect 5632 29164 5684 29170
rect 5632 29106 5684 29112
rect 4988 28552 5040 28558
rect 4988 28494 5040 28500
rect 5448 28552 5500 28558
rect 5448 28494 5500 28500
rect 5000 27538 5028 28494
rect 5540 28416 5592 28422
rect 5540 28358 5592 28364
rect 5552 27538 5580 28358
rect 9404 27872 9456 27878
rect 9404 27814 9456 27820
rect 10324 27872 10376 27878
rect 10324 27814 10376 27820
rect 9416 27538 9444 27814
rect 10336 27606 10364 27814
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 4988 27532 5040 27538
rect 4988 27474 5040 27480
rect 5540 27532 5592 27538
rect 5540 27474 5592 27480
rect 9404 27532 9456 27538
rect 9404 27474 9456 27480
rect 9496 27532 9548 27538
rect 9496 27474 9548 27480
rect 9508 26314 9536 27474
rect 8944 26308 8996 26314
rect 8944 26250 8996 26256
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 5080 21956 5132 21962
rect 5080 21898 5132 21904
rect 5092 21690 5120 21898
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 4896 21548 4948 21554
rect 4896 21490 4948 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3516 19440 3568 19446
rect 3516 19382 3568 19388
rect 3422 3496 3478 3505
rect 3422 3431 3478 3440
rect 3528 2145 3556 19382
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4908 17202 4936 21490
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5460 17746 5488 18022
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5552 17338 5580 17546
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 5460 14414 5488 17138
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5816 11280 5868 11286
rect 5816 11222 5868 11228
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3620 4865 3648 11154
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 3606 4856 3662 4865
rect 4214 4859 4522 4868
rect 3606 4791 3662 4800
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2530 4660 3470
rect 4540 2502 4660 2530
rect 3514 2136 3570 2145
rect 3514 2071 3570 2080
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect -10 0 102 800
rect 634 0 746 800
rect 1922 0 2034 800
rect 3210 0 3322 800
rect 3436 785 3464 1294
rect 4540 800 4568 2502
rect 5828 800 5856 11222
rect 6840 3534 6868 17682
rect 6932 16574 6960 23598
rect 8956 16590 8984 26250
rect 10796 23118 10824 29582
rect 12176 29170 12204 29582
rect 12164 29164 12216 29170
rect 12164 29106 12216 29112
rect 12636 28558 12664 42162
rect 20640 42158 20668 56306
rect 20904 51876 20956 51882
rect 20904 51818 20956 51824
rect 20628 42152 20680 42158
rect 20628 42094 20680 42100
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 20628 37868 20680 37874
rect 20628 37810 20680 37816
rect 20640 37262 20668 37810
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 20640 36786 20668 37198
rect 20916 37194 20944 51818
rect 22192 44872 22244 44878
rect 22192 44814 22244 44820
rect 22100 39500 22152 39506
rect 22100 39442 22152 39448
rect 21364 38344 21416 38350
rect 21364 38286 21416 38292
rect 22008 38344 22060 38350
rect 22112 38298 22140 39442
rect 22060 38292 22140 38298
rect 22008 38286 22140 38292
rect 21376 37330 21404 38286
rect 22020 38270 22140 38286
rect 21364 37324 21416 37330
rect 21364 37266 21416 37272
rect 22204 37262 22232 44814
rect 23848 40112 23900 40118
rect 23848 40054 23900 40060
rect 22284 39432 22336 39438
rect 22284 39374 22336 39380
rect 22296 38962 22324 39374
rect 22284 38956 22336 38962
rect 22284 38898 22336 38904
rect 22468 38888 22520 38894
rect 22468 38830 22520 38836
rect 22480 38554 22508 38830
rect 22468 38548 22520 38554
rect 22468 38490 22520 38496
rect 23860 38350 23888 40054
rect 24136 39030 24164 68342
rect 24860 60104 24912 60110
rect 24860 60046 24912 60052
rect 26976 60104 27028 60110
rect 26976 60046 27028 60052
rect 24872 58546 24900 60046
rect 26988 59090 27016 60046
rect 27160 59560 27212 59566
rect 27160 59502 27212 59508
rect 27172 59226 27200 59502
rect 27160 59220 27212 59226
rect 27160 59162 27212 59168
rect 26976 59084 27028 59090
rect 26976 59026 27028 59032
rect 24952 59016 25004 59022
rect 24952 58958 25004 58964
rect 24860 58540 24912 58546
rect 24860 58482 24912 58488
rect 24964 56506 24992 58958
rect 27160 58948 27212 58954
rect 27160 58890 27212 58896
rect 27172 58682 27200 58890
rect 27160 58676 27212 58682
rect 27160 58618 27212 58624
rect 24952 56500 25004 56506
rect 24952 56442 25004 56448
rect 27528 53984 27580 53990
rect 27528 53926 27580 53932
rect 27540 53650 27568 53926
rect 27528 53644 27580 53650
rect 27528 53586 27580 53592
rect 27896 53508 27948 53514
rect 27896 53450 27948 53456
rect 27908 53242 27936 53450
rect 27896 53236 27948 53242
rect 27896 53178 27948 53184
rect 27436 50312 27488 50318
rect 27436 50254 27488 50260
rect 27448 49842 27476 50254
rect 28276 49978 28304 68954
rect 28724 63912 28776 63918
rect 28724 63854 28776 63860
rect 28736 63578 28764 63854
rect 28724 63572 28776 63578
rect 28724 63514 28776 63520
rect 28264 49972 28316 49978
rect 28264 49914 28316 49920
rect 27436 49836 27488 49842
rect 27436 49778 27488 49784
rect 27620 49768 27672 49774
rect 27620 49710 27672 49716
rect 27632 49434 27660 49710
rect 27620 49428 27672 49434
rect 27620 49370 27672 49376
rect 28540 49224 28592 49230
rect 28540 49166 28592 49172
rect 28552 44878 28580 49166
rect 28540 44872 28592 44878
rect 28540 44814 28592 44820
rect 24860 42152 24912 42158
rect 24860 42094 24912 42100
rect 24872 41478 24900 42094
rect 24860 41472 24912 41478
rect 24860 41414 24912 41420
rect 26424 41472 26476 41478
rect 26424 41414 26476 41420
rect 24124 39024 24176 39030
rect 24124 38966 24176 38972
rect 23848 38344 23900 38350
rect 23848 38286 23900 38292
rect 22652 38276 22704 38282
rect 22652 38218 22704 38224
rect 22664 38010 22692 38218
rect 22652 38004 22704 38010
rect 22652 37946 22704 37952
rect 22560 37868 22612 37874
rect 22560 37810 22612 37816
rect 22192 37256 22244 37262
rect 22192 37198 22244 37204
rect 20904 37188 20956 37194
rect 20904 37130 20956 37136
rect 20628 36780 20680 36786
rect 20628 36722 20680 36728
rect 20640 36378 20668 36722
rect 20628 36372 20680 36378
rect 20628 36314 20680 36320
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 20628 30728 20680 30734
rect 20628 30670 20680 30676
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 12716 29096 12768 29102
rect 12716 29038 12768 29044
rect 12808 29096 12860 29102
rect 12808 29038 12860 29044
rect 12728 28762 12756 29038
rect 12716 28756 12768 28762
rect 12716 28698 12768 28704
rect 12624 28552 12676 28558
rect 12624 28494 12676 28500
rect 12820 27402 12848 29038
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 20640 28082 20668 30670
rect 20916 29714 20944 37130
rect 20904 29708 20956 29714
rect 20904 29650 20956 29656
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 12808 27396 12860 27402
rect 12808 27338 12860 27344
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 22204 26234 22232 37198
rect 22572 30802 22600 37810
rect 22560 30796 22612 30802
rect 22560 30738 22612 30744
rect 26436 30734 26464 41414
rect 28736 37942 28764 63514
rect 28828 59702 28856 71318
rect 28970 71318 29316 71346
rect 28970 71200 29082 71318
rect 28816 59696 28868 59702
rect 28816 59638 28868 59644
rect 29288 49910 29316 71318
rect 30258 71200 30370 72000
rect 31546 71200 31658 72000
rect 32834 71200 32946 72000
rect 34122 71200 34234 72000
rect 35410 71200 35522 72000
rect 36698 71346 36810 72000
rect 37986 71346 38098 72000
rect 36698 71318 36952 71346
rect 36698 71200 36810 71318
rect 29644 68332 29696 68338
rect 29644 68274 29696 68280
rect 29656 63442 29684 68274
rect 30300 68134 30328 71200
rect 31588 69442 31616 71200
rect 30576 69414 31616 69442
rect 30472 69284 30524 69290
rect 30472 69226 30524 69232
rect 30288 68128 30340 68134
rect 30288 68070 30340 68076
rect 30484 64666 30512 69226
rect 30472 64660 30524 64666
rect 30472 64602 30524 64608
rect 29736 64456 29788 64462
rect 29736 64398 29788 64404
rect 29748 63918 29776 64398
rect 29736 63912 29788 63918
rect 29736 63854 29788 63860
rect 29644 63436 29696 63442
rect 29644 63378 29696 63384
rect 30576 62762 30604 69414
rect 31392 69352 31444 69358
rect 31392 69294 31444 69300
rect 34060 69352 34112 69358
rect 34060 69294 34112 69300
rect 31116 68128 31168 68134
rect 31116 68070 31168 68076
rect 30932 65136 30984 65142
rect 30932 65078 30984 65084
rect 30944 64666 30972 65078
rect 30932 64660 30984 64666
rect 30932 64602 30984 64608
rect 30840 64388 30892 64394
rect 30840 64330 30892 64336
rect 30852 64122 30880 64330
rect 30840 64116 30892 64122
rect 30840 64058 30892 64064
rect 31128 64054 31156 68070
rect 31404 65618 31432 69294
rect 33140 68468 33192 68474
rect 33140 68410 33192 68416
rect 31392 65612 31444 65618
rect 31392 65554 31444 65560
rect 31404 65074 31432 65554
rect 31852 65544 31904 65550
rect 31852 65486 31904 65492
rect 31392 65068 31444 65074
rect 31392 65010 31444 65016
rect 31208 64592 31260 64598
rect 31208 64534 31260 64540
rect 31116 64048 31168 64054
rect 31116 63990 31168 63996
rect 30656 63572 30708 63578
rect 30656 63514 30708 63520
rect 30668 63374 30696 63514
rect 31220 63374 31248 64534
rect 30656 63368 30708 63374
rect 30656 63310 30708 63316
rect 31208 63368 31260 63374
rect 31208 63310 31260 63316
rect 30564 62756 30616 62762
rect 30564 62698 30616 62704
rect 29736 50312 29788 50318
rect 29736 50254 29788 50260
rect 29276 49904 29328 49910
rect 29276 49846 29328 49852
rect 29748 49842 29776 50254
rect 29736 49836 29788 49842
rect 29736 49778 29788 49784
rect 30380 49768 30432 49774
rect 30380 49710 30432 49716
rect 30392 49434 30420 49710
rect 30380 49428 30432 49434
rect 30380 49370 30432 49376
rect 28724 37936 28776 37942
rect 28724 37878 28776 37884
rect 28816 37800 28868 37806
rect 28816 37742 28868 37748
rect 26424 30728 26476 30734
rect 26424 30670 26476 30676
rect 27068 30728 27120 30734
rect 27068 30670 27120 30676
rect 27080 30258 27108 30670
rect 27068 30252 27120 30258
rect 27068 30194 27120 30200
rect 26240 27872 26292 27878
rect 26240 27814 26292 27820
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 23572 27600 23624 27606
rect 23572 27542 23624 27548
rect 23584 26246 23612 27542
rect 26252 27538 26280 27814
rect 26240 27532 26292 27538
rect 26240 27474 26292 27480
rect 27080 27402 27108 27814
rect 27068 27396 27120 27402
rect 27068 27338 27120 27344
rect 22112 26206 22232 26234
rect 23572 26240 23624 26246
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10796 22098 10824 22918
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 11624 21962 11652 23054
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 11612 21956 11664 21962
rect 11612 21898 11664 21904
rect 8944 16584 8996 16590
rect 6932 16546 7144 16574
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 7116 800 7144 16546
rect 8944 16526 8996 16532
rect 12360 3534 12388 22034
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12820 15026 12848 15438
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13004 14618 13032 14894
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 10980 800 11008 3470
rect 13556 800 13584 14894
rect 22112 14414 22140 26206
rect 23572 26182 23624 26188
rect 28828 24818 28856 37742
rect 31404 36174 31432 65010
rect 31864 64530 31892 65486
rect 33152 65006 33180 68410
rect 33140 65000 33192 65006
rect 33140 64942 33192 64948
rect 31852 64524 31904 64530
rect 31852 64466 31904 64472
rect 34072 64462 34100 69294
rect 34934 69116 35242 69125
rect 34934 69114 34940 69116
rect 34996 69114 35020 69116
rect 35076 69114 35100 69116
rect 35156 69114 35180 69116
rect 35236 69114 35242 69116
rect 34996 69062 34998 69114
rect 35178 69062 35180 69114
rect 34934 69060 34940 69062
rect 34996 69060 35020 69062
rect 35076 69060 35100 69062
rect 35156 69060 35180 69062
rect 35236 69060 35242 69062
rect 34934 69051 35242 69060
rect 34934 68028 35242 68037
rect 34934 68026 34940 68028
rect 34996 68026 35020 68028
rect 35076 68026 35100 68028
rect 35156 68026 35180 68028
rect 35236 68026 35242 68028
rect 34996 67974 34998 68026
rect 35178 67974 35180 68026
rect 34934 67972 34940 67974
rect 34996 67972 35020 67974
rect 35076 67972 35100 67974
rect 35156 67972 35180 67974
rect 35236 67972 35242 67974
rect 34934 67963 35242 67972
rect 34934 66940 35242 66949
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66875 35242 66884
rect 34934 65852 35242 65861
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65787 35242 65796
rect 34934 64764 35242 64773
rect 34934 64762 34940 64764
rect 34996 64762 35020 64764
rect 35076 64762 35100 64764
rect 35156 64762 35180 64764
rect 35236 64762 35242 64764
rect 34996 64710 34998 64762
rect 35178 64710 35180 64762
rect 34934 64708 34940 64710
rect 34996 64708 35020 64710
rect 35076 64708 35100 64710
rect 35156 64708 35180 64710
rect 35236 64708 35242 64710
rect 34934 64699 35242 64708
rect 31576 64456 31628 64462
rect 31576 64398 31628 64404
rect 34060 64456 34112 64462
rect 34060 64398 34112 64404
rect 34152 64456 34204 64462
rect 34152 64398 34204 64404
rect 31588 63986 31616 64398
rect 33232 64388 33284 64394
rect 33232 64330 33284 64336
rect 32588 64116 32640 64122
rect 32588 64058 32640 64064
rect 31576 63980 31628 63986
rect 31576 63922 31628 63928
rect 32312 63912 32364 63918
rect 32312 63854 32364 63860
rect 32324 63306 32352 63854
rect 32312 63300 32364 63306
rect 32312 63242 32364 63248
rect 32600 63238 32628 64058
rect 33244 63510 33272 64330
rect 33232 63504 33284 63510
rect 33232 63446 33284 63452
rect 33140 63368 33192 63374
rect 33140 63310 33192 63316
rect 32588 63232 32640 63238
rect 32588 63174 32640 63180
rect 32404 62824 32456 62830
rect 32404 62766 32456 62772
rect 32416 62490 32444 62766
rect 32404 62484 32456 62490
rect 32404 62426 32456 62432
rect 32600 55282 32628 63174
rect 33152 62286 33180 63310
rect 33140 62280 33192 62286
rect 33140 62222 33192 62228
rect 34164 60586 34192 64398
rect 34934 63676 35242 63685
rect 34934 63674 34940 63676
rect 34996 63674 35020 63676
rect 35076 63674 35100 63676
rect 35156 63674 35180 63676
rect 35236 63674 35242 63676
rect 34996 63622 34998 63674
rect 35178 63622 35180 63674
rect 34934 63620 34940 63622
rect 34996 63620 35020 63622
rect 35076 63620 35100 63622
rect 35156 63620 35180 63622
rect 35236 63620 35242 63622
rect 34934 63611 35242 63620
rect 34934 62588 35242 62597
rect 34934 62586 34940 62588
rect 34996 62586 35020 62588
rect 35076 62586 35100 62588
rect 35156 62586 35180 62588
rect 35236 62586 35242 62588
rect 34996 62534 34998 62586
rect 35178 62534 35180 62586
rect 34934 62532 34940 62534
rect 34996 62532 35020 62534
rect 35076 62532 35100 62534
rect 35156 62532 35180 62534
rect 35236 62532 35242 62534
rect 34934 62523 35242 62532
rect 34934 61500 35242 61509
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61435 35242 61444
rect 34152 60580 34204 60586
rect 34152 60522 34204 60528
rect 34934 60412 35242 60421
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60347 35242 60356
rect 34934 59324 35242 59333
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59259 35242 59268
rect 34934 58236 35242 58245
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58171 35242 58180
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 33048 55616 33100 55622
rect 33048 55558 33100 55564
rect 32588 55276 32640 55282
rect 32588 55218 32640 55224
rect 33060 55214 33088 55558
rect 33048 55208 33100 55214
rect 33048 55150 33100 55156
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34888 51400 34940 51406
rect 34888 51342 34940 51348
rect 34900 50930 34928 51342
rect 36728 51264 36780 51270
rect 36728 51206 36780 51212
rect 36740 50998 36768 51206
rect 36728 50992 36780 50998
rect 36728 50934 36780 50940
rect 34888 50924 34940 50930
rect 34888 50866 34940 50872
rect 35348 50856 35400 50862
rect 35348 50798 35400 50804
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 35360 50522 35388 50798
rect 35348 50516 35400 50522
rect 35348 50458 35400 50464
rect 35440 50312 35492 50318
rect 35440 50254 35492 50260
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35348 39840 35400 39846
rect 35348 39782 35400 39788
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35360 39506 35388 39782
rect 35348 39500 35400 39506
rect 35348 39442 35400 39448
rect 34888 39364 34940 39370
rect 34888 39306 34940 39312
rect 34900 39098 34928 39306
rect 34888 39092 34940 39098
rect 34888 39034 34940 39040
rect 34704 38956 34756 38962
rect 34704 38898 34756 38904
rect 32312 38344 32364 38350
rect 32312 38286 32364 38292
rect 32324 37874 32352 38286
rect 33508 38276 33560 38282
rect 33508 38218 33560 38224
rect 33520 38010 33548 38218
rect 33508 38004 33560 38010
rect 33508 37946 33560 37952
rect 32312 37868 32364 37874
rect 32312 37810 32364 37816
rect 34716 36718 34744 38898
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35452 37194 35480 50254
rect 36924 39506 36952 71318
rect 37986 71318 38608 71346
rect 37986 71200 38098 71318
rect 38580 68762 38608 71318
rect 39274 71200 39386 72000
rect 40562 71200 40674 72000
rect 41850 71200 41962 72000
rect 43138 71200 43250 72000
rect 44426 71200 44538 72000
rect 45714 71200 45826 72000
rect 47002 71482 47114 72000
rect 47002 71466 47440 71482
rect 47002 71460 47452 71466
rect 47002 71454 47400 71460
rect 47002 71200 47114 71454
rect 47400 71402 47452 71408
rect 47646 71346 47758 72000
rect 48228 71460 48280 71466
rect 48228 71402 48280 71408
rect 47228 71318 47758 71346
rect 38580 68734 38700 68762
rect 38568 68468 38620 68474
rect 38568 68410 38620 68416
rect 37924 68128 37976 68134
rect 37924 68070 37976 68076
rect 37464 66632 37516 66638
rect 37464 66574 37516 66580
rect 37476 66162 37504 66574
rect 37464 66156 37516 66162
rect 37464 66098 37516 66104
rect 37740 66088 37792 66094
rect 37740 66030 37792 66036
rect 37752 65754 37780 66030
rect 37740 65748 37792 65754
rect 37740 65690 37792 65696
rect 37936 64054 37964 68070
rect 37924 64048 37976 64054
rect 37924 63990 37976 63996
rect 38476 62144 38528 62150
rect 38476 62086 38528 62092
rect 37280 61804 37332 61810
rect 37280 61746 37332 61752
rect 37292 55282 37320 61746
rect 38488 58546 38516 62086
rect 37924 58540 37976 58546
rect 37924 58482 37976 58488
rect 38476 58540 38528 58546
rect 38476 58482 38528 58488
rect 37280 55276 37332 55282
rect 37280 55218 37332 55224
rect 37292 50402 37320 55218
rect 37292 50374 37412 50402
rect 37280 45960 37332 45966
rect 37280 45902 37332 45908
rect 37292 45490 37320 45902
rect 37280 45484 37332 45490
rect 37280 45426 37332 45432
rect 36912 39500 36964 39506
rect 36912 39442 36964 39448
rect 35440 37188 35492 37194
rect 35440 37130 35492 37136
rect 34704 36712 34756 36718
rect 34704 36654 34756 36660
rect 31392 36168 31444 36174
rect 31392 36110 31444 36116
rect 28908 30660 28960 30666
rect 28908 30602 28960 30608
rect 28816 24812 28868 24818
rect 28816 24754 28868 24760
rect 28356 24608 28408 24614
rect 28356 24550 28408 24556
rect 28540 24608 28592 24614
rect 28540 24550 28592 24556
rect 28368 23730 28396 24550
rect 28552 23798 28580 24550
rect 28540 23792 28592 23798
rect 28540 23734 28592 23740
rect 28356 23724 28408 23730
rect 28356 23666 28408 23672
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 19444 13938 19472 14350
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19628 13530 19656 13806
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 22112 13326 22140 14350
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22204 14006 22232 14214
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22204 13530 22232 13806
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19984 11076 20036 11082
rect 19984 11018 20036 11024
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14844 800 14872 2858
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 11018
rect 22572 800 22600 13806
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 11150 24624 11494
rect 26896 11150 26924 12174
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 24768 11076 24820 11082
rect 24768 11018 24820 11024
rect 24780 10962 24808 11018
rect 26240 11008 26292 11014
rect 24780 10934 24900 10962
rect 26240 10950 26292 10956
rect 24872 10810 24900 10934
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 26056 10464 26108 10470
rect 26056 10406 26108 10412
rect 26068 10130 26096 10406
rect 26252 10130 26280 10950
rect 26896 10674 26924 11086
rect 26884 10668 26936 10674
rect 26884 10610 26936 10616
rect 26056 10124 26108 10130
rect 26056 10066 26108 10072
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 27804 9988 27856 9994
rect 27804 9930 27856 9936
rect 27068 8900 27120 8906
rect 27068 8842 27120 8848
rect 27080 8634 27108 8842
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 24492 3596 24544 3602
rect 24492 3538 24544 3544
rect 24504 800 24532 3538
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26436 3058 26464 3470
rect 27068 3460 27120 3466
rect 27068 3402 27120 3408
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 26988 2446 27016 2994
rect 27080 2650 27108 3402
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 27632 2650 27660 2926
rect 27068 2644 27120 2650
rect 27068 2586 27120 2592
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 26976 2440 27028 2446
rect 26976 2382 27028 2388
rect 27816 1358 27844 9930
rect 28920 3602 28948 30602
rect 34716 25906 34744 36654
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 37096 35488 37148 35494
rect 37096 35430 37148 35436
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 37108 35154 37136 35430
rect 37096 35148 37148 35154
rect 37096 35090 37148 35096
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 37384 32502 37412 50374
rect 37464 45416 37516 45422
rect 37464 45358 37516 45364
rect 37476 45082 37504 45358
rect 37464 45076 37516 45082
rect 37464 45018 37516 45024
rect 37740 44396 37792 44402
rect 37740 44338 37792 44344
rect 37752 42158 37780 44338
rect 37936 44334 37964 58482
rect 38200 53100 38252 53106
rect 38200 53042 38252 53048
rect 38212 50318 38240 53042
rect 38200 50312 38252 50318
rect 38200 50254 38252 50260
rect 38580 45554 38608 68410
rect 38672 66094 38700 68734
rect 39316 68134 39344 71200
rect 41892 68950 41920 71200
rect 41880 68944 41932 68950
rect 41880 68886 41932 68892
rect 40684 68672 40736 68678
rect 40684 68614 40736 68620
rect 39304 68128 39356 68134
rect 39304 68070 39356 68076
rect 38660 66088 38712 66094
rect 38660 66030 38712 66036
rect 38844 53984 38896 53990
rect 38844 53926 38896 53932
rect 38856 53106 38884 53926
rect 40696 53174 40724 68614
rect 43180 67658 43208 71200
rect 44468 68406 44496 71200
rect 44456 68400 44508 68406
rect 44456 68342 44508 68348
rect 43168 67652 43220 67658
rect 43168 67594 43220 67600
rect 44180 67652 44232 67658
rect 45756 67634 45784 71200
rect 46756 69216 46808 69222
rect 46756 69158 46808 69164
rect 46572 69012 46624 69018
rect 46572 68954 46624 68960
rect 46584 68678 46612 68954
rect 46768 68882 46796 69158
rect 46756 68876 46808 68882
rect 46756 68818 46808 68824
rect 46572 68672 46624 68678
rect 46572 68614 46624 68620
rect 44180 67594 44232 67600
rect 45480 67606 45784 67634
rect 43812 66632 43864 66638
rect 43812 66574 43864 66580
rect 43824 66162 43852 66574
rect 43812 66156 43864 66162
rect 43812 66098 43864 66104
rect 43996 66088 44048 66094
rect 43996 66030 44048 66036
rect 44008 65754 44036 66030
rect 43996 65748 44048 65754
rect 43996 65690 44048 65696
rect 42616 65544 42668 65550
rect 42616 65486 42668 65492
rect 43904 65544 43956 65550
rect 43904 65486 43956 65492
rect 42628 65074 42656 65486
rect 43536 65476 43588 65482
rect 43536 65418 43588 65424
rect 42616 65068 42668 65074
rect 42616 65010 42668 65016
rect 42800 65000 42852 65006
rect 42800 64942 42852 64948
rect 42812 64666 42840 64942
rect 42800 64660 42852 64666
rect 42800 64602 42852 64608
rect 40684 53168 40736 53174
rect 40684 53110 40736 53116
rect 38844 53100 38896 53106
rect 38844 53042 38896 53048
rect 41604 49224 41656 49230
rect 41604 49166 41656 49172
rect 38488 45526 38608 45554
rect 38488 45422 38516 45526
rect 38476 45416 38528 45422
rect 38476 45358 38528 45364
rect 37924 44328 37976 44334
rect 37924 44270 37976 44276
rect 37740 42152 37792 42158
rect 37740 42094 37792 42100
rect 38844 36780 38896 36786
rect 38844 36722 38896 36728
rect 38108 36576 38160 36582
rect 38108 36518 38160 36524
rect 38120 35698 38148 36518
rect 38856 35834 38884 36722
rect 38936 36576 38988 36582
rect 38936 36518 38988 36524
rect 38844 35828 38896 35834
rect 38844 35770 38896 35776
rect 38948 35766 38976 36518
rect 38936 35760 38988 35766
rect 38936 35702 38988 35708
rect 38108 35692 38160 35698
rect 38108 35634 38160 35640
rect 39764 35624 39816 35630
rect 39764 35566 39816 35572
rect 37372 32496 37424 32502
rect 37372 32438 37424 32444
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34704 25900 34756 25906
rect 34704 25842 34756 25848
rect 34796 25696 34848 25702
rect 34796 25638 34848 25644
rect 34808 25362 34836 25638
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34796 25356 34848 25362
rect 34796 25298 34848 25304
rect 34888 25288 34940 25294
rect 34888 25230 34940 25236
rect 34900 24818 34928 25230
rect 36728 25220 36780 25226
rect 36728 25162 36780 25168
rect 34888 24812 34940 24818
rect 34888 24754 34940 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 36740 23322 36768 25162
rect 36728 23316 36780 23322
rect 36728 23258 36780 23264
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 32128 19848 32180 19854
rect 32128 19790 32180 19796
rect 32140 19378 32168 19790
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 32312 19304 32364 19310
rect 32312 19246 32364 19252
rect 32324 18970 32352 19246
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 32312 18964 32364 18970
rect 32312 18906 32364 18912
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35624 13184 35676 13190
rect 35624 13126 35676 13132
rect 35440 12640 35492 12646
rect 35440 12582 35492 12588
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35452 12306 35480 12582
rect 35636 12306 35664 13126
rect 35440 12300 35492 12306
rect 35440 12242 35492 12248
rect 35624 12300 35676 12306
rect 35624 12242 35676 12248
rect 36084 12300 36136 12306
rect 36084 12242 36136 12248
rect 34428 12096 34480 12102
rect 34428 12038 34480 12044
rect 34440 11830 34468 12038
rect 34428 11824 34480 11830
rect 34428 11766 34480 11772
rect 34796 11688 34848 11694
rect 34796 11630 34848 11636
rect 30104 11552 30156 11558
rect 30104 11494 30156 11500
rect 30116 11150 30144 11494
rect 30104 11144 30156 11150
rect 30104 11086 30156 11092
rect 30656 11076 30708 11082
rect 30656 11018 30708 11024
rect 30668 10810 30696 11018
rect 30656 10804 30708 10810
rect 30656 10746 30708 10752
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 27804 1352 27856 1358
rect 27804 1294 27856 1300
rect 34808 800 34836 11630
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35072 11076 35124 11082
rect 35072 11018 35124 11024
rect 35084 10810 35112 11018
rect 35072 10804 35124 10810
rect 35072 10746 35124 10752
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 36096 800 36124 12242
rect 39776 6914 39804 35566
rect 41616 33454 41644 49166
rect 43444 48136 43496 48142
rect 43444 48078 43496 48084
rect 43456 47666 43484 48078
rect 43444 47660 43496 47666
rect 43444 47602 43496 47608
rect 43548 47122 43576 65418
rect 43916 64462 43944 65486
rect 44192 65006 44220 67594
rect 45480 66094 45508 67606
rect 45468 66088 45520 66094
rect 45468 66030 45520 66036
rect 44180 65000 44232 65006
rect 44180 64942 44232 64948
rect 43904 64456 43956 64462
rect 43904 64398 43956 64404
rect 43628 48544 43680 48550
rect 43628 48486 43680 48492
rect 43640 47734 43668 48486
rect 43916 48278 43944 64398
rect 44180 63368 44232 63374
rect 44180 63310 44232 63316
rect 44192 61198 44220 63310
rect 46480 62688 46532 62694
rect 46480 62630 46532 62636
rect 46492 62354 46520 62630
rect 46480 62348 46532 62354
rect 46480 62290 46532 62296
rect 46664 62212 46716 62218
rect 46664 62154 46716 62160
rect 46676 61946 46704 62154
rect 46664 61940 46716 61946
rect 46664 61882 46716 61888
rect 44180 61192 44232 61198
rect 44180 61134 44232 61140
rect 44364 61192 44416 61198
rect 44364 61134 44416 61140
rect 44376 48822 44404 61134
rect 47228 60246 47256 71318
rect 47646 71200 47758 71318
rect 48240 62354 48268 71402
rect 48934 71346 49046 72000
rect 50222 71346 50334 72000
rect 48332 71318 49046 71346
rect 48228 62348 48280 62354
rect 48228 62290 48280 62296
rect 47216 60240 47268 60246
rect 47216 60182 47268 60188
rect 47676 60036 47728 60042
rect 47676 59978 47728 59984
rect 47688 59770 47716 59978
rect 47676 59764 47728 59770
rect 47676 59706 47728 59712
rect 48332 57322 48360 71318
rect 48934 71200 49046 71318
rect 49804 71318 50334 71346
rect 49148 68808 49200 68814
rect 49148 68750 49200 68756
rect 49160 68338 49188 68750
rect 49148 68332 49200 68338
rect 49148 68274 49200 68280
rect 49160 63034 49188 68274
rect 49700 63368 49752 63374
rect 49700 63310 49752 63316
rect 49148 63028 49200 63034
rect 49148 62970 49200 62976
rect 49712 62898 49740 63310
rect 49516 62892 49568 62898
rect 49516 62834 49568 62840
rect 49700 62892 49752 62898
rect 49700 62834 49752 62840
rect 48504 59628 48556 59634
rect 48504 59570 48556 59576
rect 48412 57928 48464 57934
rect 48412 57870 48464 57876
rect 48424 57458 48452 57870
rect 48412 57452 48464 57458
rect 48412 57394 48464 57400
rect 48320 57316 48372 57322
rect 48320 57258 48372 57264
rect 48516 56846 48544 59570
rect 48596 57384 48648 57390
rect 48596 57326 48648 57332
rect 48608 57050 48636 57326
rect 48596 57044 48648 57050
rect 48596 56986 48648 56992
rect 48504 56840 48556 56846
rect 48504 56782 48556 56788
rect 49056 56840 49108 56846
rect 49056 56782 49108 56788
rect 49068 55282 49096 56782
rect 49056 55276 49108 55282
rect 49056 55218 49108 55224
rect 45376 52964 45428 52970
rect 45376 52906 45428 52912
rect 44364 48816 44416 48822
rect 44364 48758 44416 48764
rect 44180 48748 44232 48754
rect 44180 48690 44232 48696
rect 43904 48272 43956 48278
rect 43904 48214 43956 48220
rect 43628 47728 43680 47734
rect 43628 47670 43680 47676
rect 43536 47116 43588 47122
rect 43536 47058 43588 47064
rect 43812 47116 43864 47122
rect 43812 47058 43864 47064
rect 43824 44402 43852 47058
rect 43812 44396 43864 44402
rect 43812 44338 43864 44344
rect 43536 42152 43588 42158
rect 43536 42094 43588 42100
rect 42340 33992 42392 33998
rect 42340 33934 42392 33940
rect 42892 33992 42944 33998
rect 42892 33934 42944 33940
rect 42352 33522 42380 33934
rect 42708 33924 42760 33930
rect 42708 33866 42760 33872
rect 42340 33516 42392 33522
rect 42340 33458 42392 33464
rect 41604 33448 41656 33454
rect 41604 33390 41656 33396
rect 41616 28082 41644 33390
rect 42352 32910 42380 33458
rect 42340 32904 42392 32910
rect 42340 32846 42392 32852
rect 42352 32434 42380 32846
rect 42340 32428 42392 32434
rect 42340 32370 42392 32376
rect 42352 30734 42380 32370
rect 42720 31822 42748 33866
rect 42904 33522 42932 33934
rect 42892 33516 42944 33522
rect 42892 33458 42944 33464
rect 43076 33448 43128 33454
rect 43076 33390 43128 33396
rect 43088 33114 43116 33390
rect 43076 33108 43128 33114
rect 43076 33050 43128 33056
rect 42984 32904 43036 32910
rect 42984 32846 43036 32852
rect 42708 31816 42760 31822
rect 42708 31758 42760 31764
rect 42616 31680 42668 31686
rect 42616 31622 42668 31628
rect 42628 31414 42656 31622
rect 42616 31408 42668 31414
rect 42616 31350 42668 31356
rect 42800 31136 42852 31142
rect 42800 31078 42852 31084
rect 42340 30728 42392 30734
rect 42340 30670 42392 30676
rect 42352 30326 42380 30670
rect 42812 30666 42840 31078
rect 42800 30660 42852 30666
rect 42800 30602 42852 30608
rect 42340 30320 42392 30326
rect 42340 30262 42392 30268
rect 42996 30054 43024 32846
rect 43352 31136 43404 31142
rect 43352 31078 43404 31084
rect 42984 30048 43036 30054
rect 42984 29990 43036 29996
rect 41604 28076 41656 28082
rect 41604 28018 41656 28024
rect 38672 6886 39804 6914
rect 38672 800 38700 6886
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 39580 2984 39632 2990
rect 39580 2926 39632 2932
rect 39948 2984 40000 2990
rect 39948 2926 40000 2932
rect 39592 2650 39620 2926
rect 39580 2644 39632 2650
rect 39580 2586 39632 2592
rect 39960 800 39988 2926
rect 40696 2650 40724 3470
rect 41788 3460 41840 3466
rect 41788 3402 41840 3408
rect 41236 3392 41288 3398
rect 41236 3334 41288 3340
rect 40684 2644 40736 2650
rect 40684 2586 40736 2592
rect 41248 800 41276 3334
rect 41800 3194 41828 3402
rect 41788 3188 41840 3194
rect 41788 3130 41840 3136
rect 42996 3058 43024 29990
rect 43364 10062 43392 31078
rect 43548 28558 43576 42094
rect 43824 32978 43852 44338
rect 43916 36786 43944 48214
rect 44192 48074 44220 48690
rect 44180 48068 44232 48074
rect 44180 48010 44232 48016
rect 44192 47122 44220 48010
rect 44180 47116 44232 47122
rect 44180 47058 44232 47064
rect 44088 44192 44140 44198
rect 44088 44134 44140 44140
rect 44100 42226 44128 44134
rect 44088 42220 44140 42226
rect 44088 42162 44140 42168
rect 44376 41138 44404 48758
rect 45284 48068 45336 48074
rect 45284 48010 45336 48016
rect 44364 41132 44416 41138
rect 44364 41074 44416 41080
rect 44376 38962 44404 41074
rect 44364 38956 44416 38962
rect 44364 38898 44416 38904
rect 45192 38752 45244 38758
rect 45192 38694 45244 38700
rect 45204 38418 45232 38694
rect 45192 38412 45244 38418
rect 45192 38354 45244 38360
rect 43904 36780 43956 36786
rect 43904 36722 43956 36728
rect 44088 33380 44140 33386
rect 44088 33322 44140 33328
rect 43812 32972 43864 32978
rect 43812 32914 43864 32920
rect 43824 32434 43852 32914
rect 44100 32910 44128 33322
rect 44088 32904 44140 32910
rect 44088 32846 44140 32852
rect 44088 32768 44140 32774
rect 44088 32710 44140 32716
rect 44100 32502 44128 32710
rect 44088 32496 44140 32502
rect 44088 32438 44140 32444
rect 43812 32428 43864 32434
rect 43812 32370 43864 32376
rect 43628 29640 43680 29646
rect 43628 29582 43680 29588
rect 43640 29170 43668 29582
rect 43628 29164 43680 29170
rect 43628 29106 43680 29112
rect 43812 29096 43864 29102
rect 43812 29038 43864 29044
rect 45192 29096 45244 29102
rect 45192 29038 45244 29044
rect 43824 28762 43852 29038
rect 43812 28756 43864 28762
rect 43812 28698 43864 28704
rect 43536 28552 43588 28558
rect 43536 28494 43588 28500
rect 43352 10056 43404 10062
rect 43352 9998 43404 10004
rect 43364 8498 43392 9998
rect 43444 9920 43496 9926
rect 43444 9862 43496 9868
rect 43456 9654 43484 9862
rect 43444 9648 43496 9654
rect 43444 9590 43496 9596
rect 43536 9512 43588 9518
rect 43536 9454 43588 9460
rect 43812 9512 43864 9518
rect 43812 9454 43864 9460
rect 43548 9178 43576 9454
rect 43536 9172 43588 9178
rect 43536 9114 43588 9120
rect 43352 8492 43404 8498
rect 43352 8434 43404 8440
rect 41696 3052 41748 3058
rect 41696 2994 41748 3000
rect 42984 3052 43036 3058
rect 42984 2994 43036 3000
rect 41708 2446 41736 2994
rect 41696 2440 41748 2446
rect 41696 2382 41748 2388
rect 43824 800 43852 9454
rect 45204 4146 45232 29038
rect 45296 12374 45324 48010
rect 45388 47122 45416 52906
rect 45560 51400 45612 51406
rect 45560 51342 45612 51348
rect 45572 50998 45600 51342
rect 45560 50992 45612 50998
rect 45560 50934 45612 50940
rect 45560 50856 45612 50862
rect 45560 50798 45612 50804
rect 45572 50522 45600 50798
rect 45560 50516 45612 50522
rect 45560 50458 45612 50464
rect 47584 50312 47636 50318
rect 47584 50254 47636 50260
rect 45376 47116 45428 47122
rect 45376 47058 45428 47064
rect 45388 18766 45416 47058
rect 47596 45354 47624 50254
rect 48780 45484 48832 45490
rect 48780 45426 48832 45432
rect 47584 45348 47636 45354
rect 47584 45290 47636 45296
rect 48792 44198 48820 45426
rect 48780 44192 48832 44198
rect 48780 44134 48832 44140
rect 48792 39030 48820 44134
rect 48780 39024 48832 39030
rect 48780 38966 48832 38972
rect 46388 38888 46440 38894
rect 46388 38830 46440 38836
rect 46400 37874 46428 38830
rect 46848 38276 46900 38282
rect 46848 38218 46900 38224
rect 46388 37868 46440 37874
rect 46388 37810 46440 37816
rect 45468 32360 45520 32366
rect 45468 32302 45520 32308
rect 45376 18760 45428 18766
rect 45376 18702 45428 18708
rect 45284 12368 45336 12374
rect 45284 12310 45336 12316
rect 45192 4140 45244 4146
rect 45192 4082 45244 4088
rect 45100 4072 45152 4078
rect 45100 4014 45152 4020
rect 45112 800 45140 4014
rect 45480 3466 45508 32302
rect 46860 4078 46888 38218
rect 48792 37874 48820 38966
rect 48780 37868 48832 37874
rect 48780 37810 48832 37816
rect 48964 37800 49016 37806
rect 48964 37742 49016 37748
rect 47584 32292 47636 32298
rect 47584 32234 47636 32240
rect 47596 22642 47624 32234
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 48976 10674 49004 37742
rect 49068 33930 49096 55218
rect 49528 45490 49556 62834
rect 49804 62762 49832 71318
rect 50222 71200 50334 71318
rect 51510 71200 51622 72000
rect 52798 71200 52910 72000
rect 54086 71200 54198 72000
rect 55374 71200 55486 72000
rect 56662 71200 56774 72000
rect 57950 71200 58062 72000
rect 59238 71200 59350 72000
rect 60526 71200 60638 72000
rect 61814 71200 61926 72000
rect 63102 71200 63214 72000
rect 64390 71200 64502 72000
rect 65678 71346 65790 72000
rect 65352 71318 65790 71346
rect 50294 69660 50602 69669
rect 50294 69658 50300 69660
rect 50356 69658 50380 69660
rect 50436 69658 50460 69660
rect 50516 69658 50540 69660
rect 50596 69658 50602 69660
rect 50356 69606 50358 69658
rect 50538 69606 50540 69658
rect 50294 69604 50300 69606
rect 50356 69604 50380 69606
rect 50436 69604 50460 69606
rect 50516 69604 50540 69606
rect 50596 69604 50602 69606
rect 50294 69595 50602 69604
rect 51264 69216 51316 69222
rect 51264 69158 51316 69164
rect 51276 68882 51304 69158
rect 51552 68882 51580 71200
rect 52840 69018 52868 71200
rect 52828 69012 52880 69018
rect 52828 68954 52880 68960
rect 51264 68876 51316 68882
rect 51264 68818 51316 68824
rect 51540 68876 51592 68882
rect 51540 68818 51592 68824
rect 51172 68740 51224 68746
rect 51172 68682 51224 68688
rect 50294 68572 50602 68581
rect 50294 68570 50300 68572
rect 50356 68570 50380 68572
rect 50436 68570 50460 68572
rect 50516 68570 50540 68572
rect 50596 68570 50602 68572
rect 50356 68518 50358 68570
rect 50538 68518 50540 68570
rect 50294 68516 50300 68518
rect 50356 68516 50380 68518
rect 50436 68516 50460 68518
rect 50516 68516 50540 68518
rect 50596 68516 50602 68518
rect 50294 68507 50602 68516
rect 51184 68474 51212 68682
rect 53288 68672 53340 68678
rect 53288 68614 53340 68620
rect 51172 68468 51224 68474
rect 51172 68410 51224 68416
rect 50294 67484 50602 67493
rect 50294 67482 50300 67484
rect 50356 67482 50380 67484
rect 50436 67482 50460 67484
rect 50516 67482 50540 67484
rect 50596 67482 50602 67484
rect 50356 67430 50358 67482
rect 50538 67430 50540 67482
rect 50294 67428 50300 67430
rect 50356 67428 50380 67430
rect 50436 67428 50460 67430
rect 50516 67428 50540 67430
rect 50596 67428 50602 67430
rect 50294 67419 50602 67428
rect 50294 66396 50602 66405
rect 50294 66394 50300 66396
rect 50356 66394 50380 66396
rect 50436 66394 50460 66396
rect 50516 66394 50540 66396
rect 50596 66394 50602 66396
rect 50356 66342 50358 66394
rect 50538 66342 50540 66394
rect 50294 66340 50300 66342
rect 50356 66340 50380 66342
rect 50436 66340 50460 66342
rect 50516 66340 50540 66342
rect 50596 66340 50602 66342
rect 50294 66331 50602 66340
rect 50294 65308 50602 65317
rect 50294 65306 50300 65308
rect 50356 65306 50380 65308
rect 50436 65306 50460 65308
rect 50516 65306 50540 65308
rect 50596 65306 50602 65308
rect 50356 65254 50358 65306
rect 50538 65254 50540 65306
rect 50294 65252 50300 65254
rect 50356 65252 50380 65254
rect 50436 65252 50460 65254
rect 50516 65252 50540 65254
rect 50596 65252 50602 65254
rect 50294 65243 50602 65252
rect 50294 64220 50602 64229
rect 50294 64218 50300 64220
rect 50356 64218 50380 64220
rect 50436 64218 50460 64220
rect 50516 64218 50540 64220
rect 50596 64218 50602 64220
rect 50356 64166 50358 64218
rect 50538 64166 50540 64218
rect 50294 64164 50300 64166
rect 50356 64164 50380 64166
rect 50436 64164 50460 64166
rect 50516 64164 50540 64166
rect 50596 64164 50602 64166
rect 50294 64155 50602 64164
rect 50294 63132 50602 63141
rect 50294 63130 50300 63132
rect 50356 63130 50380 63132
rect 50436 63130 50460 63132
rect 50516 63130 50540 63132
rect 50596 63130 50602 63132
rect 50356 63078 50358 63130
rect 50538 63078 50540 63130
rect 50294 63076 50300 63078
rect 50356 63076 50380 63078
rect 50436 63076 50460 63078
rect 50516 63076 50540 63078
rect 50596 63076 50602 63078
rect 50294 63067 50602 63076
rect 50252 62824 50304 62830
rect 50252 62766 50304 62772
rect 49792 62756 49844 62762
rect 49792 62698 49844 62704
rect 50264 62490 50292 62766
rect 50252 62484 50304 62490
rect 50252 62426 50304 62432
rect 50294 62044 50602 62053
rect 50294 62042 50300 62044
rect 50356 62042 50380 62044
rect 50436 62042 50460 62044
rect 50516 62042 50540 62044
rect 50596 62042 50602 62044
rect 50356 61990 50358 62042
rect 50538 61990 50540 62042
rect 50294 61988 50300 61990
rect 50356 61988 50380 61990
rect 50436 61988 50460 61990
rect 50516 61988 50540 61990
rect 50596 61988 50602 61990
rect 50294 61979 50602 61988
rect 50294 60956 50602 60965
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60891 50602 60900
rect 50294 59868 50602 59877
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59803 50602 59812
rect 50294 58780 50602 58789
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58715 50602 58724
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 51448 53984 51500 53990
rect 51448 53926 51500 53932
rect 51460 53650 51488 53926
rect 51448 53644 51500 53650
rect 51448 53586 51500 53592
rect 51356 53508 51408 53514
rect 51356 53450 51408 53456
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 51368 53242 51396 53450
rect 51356 53236 51408 53242
rect 51356 53178 51408 53184
rect 51080 53100 51132 53106
rect 51080 53042 51132 53048
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 49516 45484 49568 45490
rect 49516 45426 49568 45432
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 49056 33924 49108 33930
rect 49056 33866 49108 33872
rect 49068 31346 49096 33866
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 51092 33114 51120 53042
rect 51356 51808 51408 51814
rect 51356 51750 51408 51756
rect 51368 51474 51396 51750
rect 53300 51474 53328 68614
rect 54128 68474 54156 71200
rect 55416 69426 55444 71200
rect 55404 69420 55456 69426
rect 55404 69362 55456 69368
rect 56704 68950 56732 71200
rect 57992 69306 58020 71200
rect 57992 69278 59124 69306
rect 56968 69216 57020 69222
rect 56968 69158 57020 69164
rect 58992 69216 59044 69222
rect 58992 69158 59044 69164
rect 56692 68944 56744 68950
rect 56692 68886 56744 68892
rect 56980 68882 57008 69158
rect 56968 68876 57020 68882
rect 56968 68818 57020 68824
rect 58900 68808 58952 68814
rect 58900 68750 58952 68756
rect 56416 68740 56468 68746
rect 56416 68682 56468 68688
rect 56428 68474 56456 68682
rect 54116 68468 54168 68474
rect 54116 68410 54168 68416
rect 56416 68468 56468 68474
rect 56416 68410 56468 68416
rect 53380 68400 53432 68406
rect 53380 68342 53432 68348
rect 51356 51468 51408 51474
rect 51356 51410 51408 51416
rect 53288 51468 53340 51474
rect 53288 51410 53340 51416
rect 51540 51332 51592 51338
rect 51540 51274 51592 51280
rect 51552 51066 51580 51274
rect 51540 51060 51592 51066
rect 51540 51002 51592 51008
rect 53196 50924 53248 50930
rect 53196 50866 53248 50872
rect 53208 48754 53236 50866
rect 53196 48748 53248 48754
rect 53196 48690 53248 48696
rect 53208 48074 53236 48690
rect 53196 48068 53248 48074
rect 53196 48010 53248 48016
rect 52092 44328 52144 44334
rect 52092 44270 52144 44276
rect 52104 43790 52132 44270
rect 52092 43784 52144 43790
rect 52092 43726 52144 43732
rect 52736 43784 52788 43790
rect 52736 43726 52788 43732
rect 52104 42702 52132 43726
rect 52748 43314 52776 43726
rect 52736 43308 52788 43314
rect 52736 43250 52788 43256
rect 52092 42696 52144 42702
rect 52092 42638 52144 42644
rect 51540 38344 51592 38350
rect 51540 38286 51592 38292
rect 51172 37868 51224 37874
rect 51172 37810 51224 37816
rect 51080 33108 51132 33114
rect 51080 33050 51132 33056
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 49056 31340 49108 31346
rect 49056 31282 49108 31288
rect 51184 31142 51212 37810
rect 51264 37664 51316 37670
rect 51264 37606 51316 37612
rect 51276 37194 51304 37606
rect 51552 37330 51580 38286
rect 51540 37324 51592 37330
rect 51540 37266 51592 37272
rect 53392 37262 53420 68342
rect 58912 68270 58940 68750
rect 59004 68338 59032 69158
rect 58992 68332 59044 68338
rect 58992 68274 59044 68280
rect 58900 68264 58952 68270
rect 58900 68206 58952 68212
rect 58624 68128 58676 68134
rect 58624 68070 58676 68076
rect 55956 64864 56008 64870
rect 55956 64806 56008 64812
rect 55968 64530 55996 64806
rect 55956 64524 56008 64530
rect 55956 64466 56008 64472
rect 55864 64388 55916 64394
rect 55864 64330 55916 64336
rect 55876 64122 55904 64330
rect 55864 64116 55916 64122
rect 55864 64058 55916 64064
rect 55588 63980 55640 63986
rect 55588 63922 55640 63928
rect 54484 62280 54536 62286
rect 54484 62222 54536 62228
rect 54496 61810 54524 62222
rect 55600 61878 55628 63922
rect 58072 63776 58124 63782
rect 58072 63718 58124 63724
rect 58084 63442 58112 63718
rect 58072 63436 58124 63442
rect 58072 63378 58124 63384
rect 57980 63300 58032 63306
rect 57980 63242 58032 63248
rect 57992 63034 58020 63242
rect 57980 63028 58032 63034
rect 57980 62970 58032 62976
rect 55588 61872 55640 61878
rect 55588 61814 55640 61820
rect 54484 61804 54536 61810
rect 54484 61746 54536 61752
rect 54668 61736 54720 61742
rect 54668 61678 54720 61684
rect 54680 61402 54708 61678
rect 54668 61396 54720 61402
rect 54668 61338 54720 61344
rect 57888 55752 57940 55758
rect 57888 55694 57940 55700
rect 57900 55282 57928 55694
rect 57888 55276 57940 55282
rect 57888 55218 57940 55224
rect 58636 53514 58664 68070
rect 58912 67250 58940 68206
rect 58900 67244 58952 67250
rect 58900 67186 58952 67192
rect 59096 63442 59124 69278
rect 59176 68672 59228 68678
rect 59176 68614 59228 68620
rect 59188 68270 59216 68614
rect 59176 68264 59228 68270
rect 59176 68206 59228 68212
rect 60568 68134 60596 71200
rect 60556 68128 60608 68134
rect 60556 68070 60608 68076
rect 60924 67720 60976 67726
rect 60924 67662 60976 67668
rect 60936 67250 60964 67662
rect 61108 67652 61160 67658
rect 61108 67594 61160 67600
rect 61120 67386 61148 67594
rect 61108 67380 61160 67386
rect 61108 67322 61160 67328
rect 60924 67244 60976 67250
rect 60924 67186 60976 67192
rect 61856 64874 61884 71200
rect 63144 68746 63172 71200
rect 64144 69012 64196 69018
rect 64144 68954 64196 68960
rect 63132 68740 63184 68746
rect 63132 68682 63184 68688
rect 62764 67652 62816 67658
rect 62764 67594 62816 67600
rect 62776 67046 62804 67594
rect 62764 67040 62816 67046
rect 62764 66982 62816 66988
rect 61856 64846 62068 64874
rect 59084 63436 59136 63442
rect 59084 63378 59136 63384
rect 58624 53508 58676 53514
rect 58624 53450 58676 53456
rect 53840 49224 53892 49230
rect 53840 49166 53892 49172
rect 53852 48754 53880 49166
rect 53840 48748 53892 48754
rect 53840 48690 53892 48696
rect 54944 42560 54996 42566
rect 54944 42502 54996 42508
rect 54956 42294 54984 42502
rect 54944 42288 54996 42294
rect 54944 42230 54996 42236
rect 56508 42152 56560 42158
rect 56508 42094 56560 42100
rect 53380 37256 53432 37262
rect 53380 37198 53432 37204
rect 51264 37188 51316 37194
rect 51264 37130 51316 37136
rect 54208 33108 54260 33114
rect 54208 33050 54260 33056
rect 51172 31136 51224 31142
rect 51172 31078 51224 31084
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 54220 28558 54248 33050
rect 54208 28552 54260 28558
rect 54208 28494 54260 28500
rect 54760 28552 54812 28558
rect 54760 28494 54812 28500
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 54772 28082 54800 28494
rect 54760 28076 54812 28082
rect 54760 28018 54812 28024
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50528 22432 50580 22438
rect 50528 22374 50580 22380
rect 51356 22432 51408 22438
rect 51356 22374 51408 22380
rect 50540 22098 50568 22374
rect 50528 22092 50580 22098
rect 50528 22034 50580 22040
rect 50804 22092 50856 22098
rect 50804 22034 50856 22040
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50816 20806 50844 22034
rect 51368 21962 51396 22374
rect 51356 21956 51408 21962
rect 51356 21898 51408 21904
rect 49792 20800 49844 20806
rect 49792 20742 49844 20748
rect 50804 20800 50856 20806
rect 50804 20742 50856 20748
rect 49804 16574 49832 20742
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 49804 16546 50936 16574
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 48964 10668 49016 10674
rect 48964 10610 49016 10616
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 47032 4140 47084 4146
rect 47032 4082 47084 4088
rect 46848 4072 46900 4078
rect 46848 4014 46900 4020
rect 45468 3460 45520 3466
rect 45468 3402 45520 3408
rect 47044 800 47072 4082
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50908 800 50936 16546
rect 54392 10056 54444 10062
rect 54392 9998 54444 10004
rect 54404 8974 54432 9998
rect 54392 8968 54444 8974
rect 54392 8910 54444 8916
rect 54760 8968 54812 8974
rect 54760 8910 54812 8916
rect 54772 8498 54800 8910
rect 54944 8832 54996 8838
rect 54944 8774 54996 8780
rect 54956 8566 54984 8774
rect 54944 8560 54996 8566
rect 54944 8502 54996 8508
rect 54760 8492 54812 8498
rect 54760 8434 54812 8440
rect 56520 3194 56548 42094
rect 57888 41064 57940 41070
rect 57888 41006 57940 41012
rect 57900 40730 57928 41006
rect 57888 40724 57940 40730
rect 57888 40666 57940 40672
rect 60464 39840 60516 39846
rect 60464 39782 60516 39788
rect 60476 39506 60504 39782
rect 62040 39506 62068 64846
rect 64156 64530 64184 68954
rect 65352 68406 65380 71318
rect 65678 71200 65790 71318
rect 66966 71200 67078 72000
rect 68254 71200 68366 72000
rect 69542 71346 69654 72000
rect 69216 71318 69654 71346
rect 65654 69116 65962 69125
rect 65654 69114 65660 69116
rect 65716 69114 65740 69116
rect 65796 69114 65820 69116
rect 65876 69114 65900 69116
rect 65956 69114 65962 69116
rect 65716 69062 65718 69114
rect 65898 69062 65900 69114
rect 65654 69060 65660 69062
rect 65716 69060 65740 69062
rect 65796 69060 65820 69062
rect 65876 69060 65900 69062
rect 65956 69060 65962 69062
rect 65654 69051 65962 69060
rect 67008 69018 67036 71200
rect 67454 70136 67510 70145
rect 67454 70071 67510 70080
rect 67468 69494 67496 70071
rect 67456 69488 67508 69494
rect 67456 69430 67508 69436
rect 66996 69012 67048 69018
rect 66996 68954 67048 68960
rect 65340 68400 65392 68406
rect 65340 68342 65392 68348
rect 68296 68270 68324 71200
rect 68284 68264 68336 68270
rect 68284 68206 68336 68212
rect 69216 68134 69244 71318
rect 69542 71200 69654 71318
rect 67732 68128 67784 68134
rect 67732 68070 67784 68076
rect 69204 68128 69256 68134
rect 69204 68070 69256 68076
rect 65654 68028 65962 68037
rect 65654 68026 65660 68028
rect 65716 68026 65740 68028
rect 65796 68026 65820 68028
rect 65876 68026 65900 68028
rect 65956 68026 65962 68028
rect 65716 67974 65718 68026
rect 65898 67974 65900 68026
rect 65654 67972 65660 67974
rect 65716 67972 65740 67974
rect 65796 67972 65820 67974
rect 65876 67972 65900 67974
rect 65956 67972 65962 67974
rect 65654 67963 65962 67972
rect 66166 67416 66222 67425
rect 66166 67351 66222 67360
rect 66180 67046 66208 67351
rect 66168 67040 66220 67046
rect 66168 66982 66220 66988
rect 65654 66940 65962 66949
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66875 65962 66884
rect 66166 66056 66222 66065
rect 66166 65991 66222 66000
rect 65654 65852 65962 65861
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65787 65962 65796
rect 65654 64764 65962 64773
rect 65654 64762 65660 64764
rect 65716 64762 65740 64764
rect 65796 64762 65820 64764
rect 65876 64762 65900 64764
rect 65956 64762 65962 64764
rect 65716 64710 65718 64762
rect 65898 64710 65900 64762
rect 65654 64708 65660 64710
rect 65716 64708 65740 64710
rect 65796 64708 65820 64710
rect 65876 64708 65900 64710
rect 65956 64708 65962 64710
rect 65654 64699 65962 64708
rect 64144 64524 64196 64530
rect 64144 64466 64196 64472
rect 65654 63676 65962 63685
rect 65654 63674 65660 63676
rect 65716 63674 65740 63676
rect 65796 63674 65820 63676
rect 65876 63674 65900 63676
rect 65956 63674 65962 63676
rect 65716 63622 65718 63674
rect 65898 63622 65900 63674
rect 65654 63620 65660 63622
rect 65716 63620 65740 63622
rect 65796 63620 65820 63622
rect 65876 63620 65900 63622
rect 65956 63620 65962 63622
rect 65654 63611 65962 63620
rect 64512 62892 64564 62898
rect 64512 62834 64564 62840
rect 64524 61810 64552 62834
rect 65156 62756 65208 62762
rect 65156 62698 65208 62704
rect 65168 61810 65196 62698
rect 65340 62688 65392 62694
rect 65340 62630 65392 62636
rect 65352 61878 65380 62630
rect 65654 62588 65962 62597
rect 65654 62586 65660 62588
rect 65716 62586 65740 62588
rect 65796 62586 65820 62588
rect 65876 62586 65900 62588
rect 65956 62586 65962 62588
rect 65716 62534 65718 62586
rect 65898 62534 65900 62586
rect 65654 62532 65660 62534
rect 65716 62532 65740 62534
rect 65796 62532 65820 62534
rect 65876 62532 65900 62534
rect 65956 62532 65962 62534
rect 65654 62523 65962 62532
rect 65800 62212 65852 62218
rect 65800 62154 65852 62160
rect 65812 61946 65840 62154
rect 66074 61976 66130 61985
rect 65800 61940 65852 61946
rect 66074 61911 66130 61920
rect 65800 61882 65852 61888
rect 65340 61872 65392 61878
rect 65340 61814 65392 61820
rect 64512 61804 64564 61810
rect 64512 61746 64564 61752
rect 65156 61804 65208 61810
rect 65156 61746 65208 61752
rect 63224 50720 63276 50726
rect 63224 50662 63276 50668
rect 63236 50386 63264 50662
rect 63224 50380 63276 50386
rect 63224 50322 63276 50328
rect 63408 50244 63460 50250
rect 63408 50186 63460 50192
rect 63420 49978 63448 50186
rect 63408 49972 63460 49978
rect 63408 49914 63460 49920
rect 62948 49836 63000 49842
rect 62948 49778 63000 49784
rect 62960 46986 62988 49778
rect 64524 48618 64552 61746
rect 66088 61742 66116 61911
rect 66076 61736 66128 61742
rect 66076 61678 66128 61684
rect 65654 61500 65962 61509
rect 65654 61498 65660 61500
rect 65716 61498 65740 61500
rect 65796 61498 65820 61500
rect 65876 61498 65900 61500
rect 65956 61498 65962 61500
rect 65716 61446 65718 61498
rect 65898 61446 65900 61498
rect 65654 61444 65660 61446
rect 65716 61444 65740 61446
rect 65796 61444 65820 61446
rect 65876 61444 65900 61446
rect 65956 61444 65962 61446
rect 65654 61435 65962 61444
rect 66074 60616 66130 60625
rect 66074 60551 66130 60560
rect 65654 60412 65962 60421
rect 65654 60410 65660 60412
rect 65716 60410 65740 60412
rect 65796 60410 65820 60412
rect 65876 60410 65900 60412
rect 65956 60410 65962 60412
rect 65716 60358 65718 60410
rect 65898 60358 65900 60410
rect 65654 60356 65660 60358
rect 65716 60356 65740 60358
rect 65796 60356 65820 60358
rect 65876 60356 65900 60358
rect 65956 60356 65962 60358
rect 65654 60347 65962 60356
rect 66088 59537 66116 60551
rect 64786 59528 64842 59537
rect 64786 59463 64842 59472
rect 66074 59528 66130 59537
rect 66074 59463 66130 59472
rect 64694 56672 64750 56681
rect 64694 56607 64750 56616
rect 64708 48822 64736 56607
rect 64800 50386 64828 59463
rect 65654 59324 65962 59333
rect 65654 59322 65660 59324
rect 65716 59322 65740 59324
rect 65796 59322 65820 59324
rect 65876 59322 65900 59324
rect 65956 59322 65962 59324
rect 65716 59270 65718 59322
rect 65898 59270 65900 59322
rect 65654 59268 65660 59270
rect 65716 59268 65740 59270
rect 65796 59268 65820 59270
rect 65876 59268 65900 59270
rect 65956 59268 65962 59270
rect 65654 59259 65962 59268
rect 65654 58236 65962 58245
rect 65654 58234 65660 58236
rect 65716 58234 65740 58236
rect 65796 58234 65820 58236
rect 65876 58234 65900 58236
rect 65956 58234 65962 58236
rect 65716 58182 65718 58234
rect 65898 58182 65900 58234
rect 65654 58180 65660 58182
rect 65716 58180 65740 58182
rect 65796 58180 65820 58182
rect 65876 58180 65900 58182
rect 65956 58180 65962 58182
rect 65654 58171 65962 58180
rect 66074 57896 66130 57905
rect 66074 57831 66130 57840
rect 65654 57148 65962 57157
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57083 65962 57092
rect 66088 56681 66116 57831
rect 66074 56672 66130 56681
rect 66074 56607 66130 56616
rect 65654 56060 65962 56069
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55995 65962 56004
rect 66076 55208 66128 55214
rect 66074 55176 66076 55185
rect 66128 55176 66130 55185
rect 66074 55111 66130 55120
rect 65654 54972 65962 54981
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54907 65962 54916
rect 65654 53884 65962 53893
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53819 65962 53828
rect 66180 53718 66208 65991
rect 67454 63336 67510 63345
rect 67454 63271 67510 63280
rect 67468 62354 67496 63271
rect 67456 62348 67508 62354
rect 67456 62290 67508 62296
rect 67744 61878 67772 68070
rect 67732 61872 67784 61878
rect 67732 61814 67784 61820
rect 66260 53984 66312 53990
rect 66260 53926 66312 53932
rect 66168 53712 66220 53718
rect 66168 53654 66220 53660
rect 66272 53650 66300 53926
rect 66260 53644 66312 53650
rect 66260 53586 66312 53592
rect 66444 53508 66496 53514
rect 66444 53450 66496 53456
rect 66456 53242 66484 53450
rect 66444 53236 66496 53242
rect 66444 53178 66496 53184
rect 67456 53100 67508 53106
rect 67456 53042 67508 53048
rect 65654 52796 65962 52805
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52731 65962 52740
rect 65654 51708 65962 51717
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51643 65962 51652
rect 66076 51264 66128 51270
rect 66076 51206 66128 51212
rect 66088 51105 66116 51206
rect 66074 51096 66130 51105
rect 66074 51031 66130 51040
rect 65654 50620 65962 50629
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50555 65962 50564
rect 64788 50380 64840 50386
rect 64788 50322 64840 50328
rect 65522 49736 65578 49745
rect 65522 49671 65578 49680
rect 64696 48816 64748 48822
rect 64696 48758 64748 48764
rect 64512 48612 64564 48618
rect 64512 48554 64564 48560
rect 64696 48612 64748 48618
rect 64696 48554 64748 48560
rect 64708 47666 64736 48554
rect 64696 47660 64748 47666
rect 64696 47602 64748 47608
rect 65340 47592 65392 47598
rect 65340 47534 65392 47540
rect 65352 47258 65380 47534
rect 65340 47252 65392 47258
rect 65340 47194 65392 47200
rect 62948 46980 63000 46986
rect 62948 46922 63000 46928
rect 60464 39500 60516 39506
rect 60464 39442 60516 39448
rect 62028 39500 62080 39506
rect 62028 39442 62080 39448
rect 60648 39364 60700 39370
rect 60648 39306 60700 39312
rect 60660 39098 60688 39306
rect 60648 39092 60700 39098
rect 60648 39034 60700 39040
rect 61844 38956 61896 38962
rect 61844 38898 61896 38904
rect 61856 32434 61884 38898
rect 62396 33312 62448 33318
rect 62396 33254 62448 33260
rect 62408 32978 62436 33254
rect 62396 32972 62448 32978
rect 62396 32914 62448 32920
rect 61936 32836 61988 32842
rect 61936 32778 61988 32784
rect 61948 32570 61976 32778
rect 61936 32564 61988 32570
rect 61936 32506 61988 32512
rect 60740 32428 60792 32434
rect 60740 32370 60792 32376
rect 61844 32428 61896 32434
rect 61844 32370 61896 32376
rect 59820 31272 59872 31278
rect 59820 31214 59872 31220
rect 59832 30938 59860 31214
rect 59820 30932 59872 30938
rect 59820 30874 59872 30880
rect 58164 24200 58216 24206
rect 58164 24142 58216 24148
rect 58176 23730 58204 24142
rect 58164 23724 58216 23730
rect 58164 23666 58216 23672
rect 58348 23656 58400 23662
rect 58348 23598 58400 23604
rect 58360 23322 58388 23598
rect 58348 23316 58400 23322
rect 58348 23258 58400 23264
rect 60752 23118 60780 32370
rect 57888 23112 57940 23118
rect 57888 23054 57940 23060
rect 60740 23112 60792 23118
rect 60740 23054 60792 23060
rect 57900 22642 57928 23054
rect 60648 23044 60700 23050
rect 60648 22986 60700 22992
rect 60660 22642 60688 22986
rect 60832 22976 60884 22982
rect 60832 22918 60884 22924
rect 60844 22710 60872 22918
rect 60832 22704 60884 22710
rect 60832 22646 60884 22652
rect 57888 22636 57940 22642
rect 57888 22578 57940 22584
rect 60648 22636 60700 22642
rect 60648 22578 60700 22584
rect 62488 22568 62540 22574
rect 62488 22510 62540 22516
rect 62500 15162 62528 22510
rect 62960 22030 62988 46922
rect 64878 42256 64934 42265
rect 64878 42191 64934 42200
rect 64892 41426 64920 42191
rect 64800 41398 64920 41426
rect 63224 39840 63276 39846
rect 63224 39782 63276 39788
rect 63236 39506 63264 39782
rect 64800 39506 64828 41398
rect 63224 39500 63276 39506
rect 63224 39442 63276 39448
rect 64788 39500 64840 39506
rect 64788 39442 64840 39448
rect 63500 39364 63552 39370
rect 63500 39306 63552 39312
rect 63512 39098 63540 39306
rect 63500 39092 63552 39098
rect 63500 39034 63552 39040
rect 63408 38956 63460 38962
rect 63408 38898 63460 38904
rect 63420 37806 63448 38898
rect 63408 37800 63460 37806
rect 63408 37742 63460 37748
rect 63420 37482 63448 37742
rect 63420 37454 63724 37482
rect 63040 35624 63092 35630
rect 63040 35566 63092 35572
rect 63052 35290 63080 35566
rect 63040 35284 63092 35290
rect 63040 35226 63092 35232
rect 63696 35086 63724 37454
rect 63776 35624 63828 35630
rect 63776 35566 63828 35572
rect 63788 35290 63816 35566
rect 63776 35284 63828 35290
rect 63776 35226 63828 35232
rect 63684 35080 63736 35086
rect 63684 35022 63736 35028
rect 63132 31272 63184 31278
rect 63132 31214 63184 31220
rect 63144 30190 63172 31214
rect 63132 30184 63184 30190
rect 63132 30126 63184 30132
rect 62948 22024 63000 22030
rect 62948 21966 63000 21972
rect 62960 17678 62988 21966
rect 63316 21888 63368 21894
rect 63316 21830 63368 21836
rect 63328 21622 63356 21830
rect 63316 21616 63368 21622
rect 63316 21558 63368 21564
rect 63132 21480 63184 21486
rect 63132 21422 63184 21428
rect 63144 21146 63172 21422
rect 63132 21140 63184 21146
rect 63132 21082 63184 21088
rect 62948 17672 63000 17678
rect 62948 17614 63000 17620
rect 63040 17672 63092 17678
rect 63040 17614 63092 17620
rect 63052 17202 63080 17614
rect 63224 17536 63276 17542
rect 63224 17478 63276 17484
rect 63236 17270 63264 17478
rect 63224 17264 63276 17270
rect 63224 17206 63276 17212
rect 63040 17196 63092 17202
rect 63040 17138 63092 17144
rect 62488 15156 62540 15162
rect 62488 15098 62540 15104
rect 63408 12232 63460 12238
rect 63408 12174 63460 12180
rect 63420 11762 63448 12174
rect 63408 11756 63460 11762
rect 63408 11698 63460 11704
rect 63316 11688 63368 11694
rect 63316 11630 63368 11636
rect 63328 11354 63356 11630
rect 63316 11348 63368 11354
rect 63316 11290 63368 11296
rect 63696 11150 63724 35022
rect 65536 33454 65564 49671
rect 65654 49532 65962 49541
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49467 65962 49476
rect 65654 48444 65962 48453
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48379 65962 48388
rect 67180 47592 67232 47598
rect 67180 47534 67232 47540
rect 65654 47356 65962 47365
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47291 65962 47300
rect 67192 46345 67220 47534
rect 67178 46336 67234 46345
rect 65654 46268 65962 46277
rect 67178 46271 67234 46280
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46203 65962 46212
rect 67468 45354 67496 53042
rect 67456 45348 67508 45354
rect 67456 45290 67508 45296
rect 66260 45280 66312 45286
rect 66260 45222 66312 45228
rect 65654 45180 65962 45189
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45115 65962 45124
rect 66272 44946 66300 45222
rect 66260 44940 66312 44946
rect 66260 44882 66312 44888
rect 66444 44804 66496 44810
rect 66444 44746 66496 44752
rect 66456 44538 66484 44746
rect 66444 44532 66496 44538
rect 66444 44474 66496 44480
rect 67468 44402 67496 45290
rect 68098 44976 68154 44985
rect 68098 44911 68100 44920
rect 68152 44911 68154 44920
rect 68100 44882 68152 44888
rect 67456 44396 67508 44402
rect 67456 44338 67508 44344
rect 65654 44092 65962 44101
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44027 65962 44036
rect 66168 43716 66220 43722
rect 66168 43658 66220 43664
rect 66180 43625 66208 43658
rect 66166 43616 66222 43625
rect 66166 43551 66222 43560
rect 65654 43004 65962 43013
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42939 65962 42948
rect 65654 41916 65962 41925
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41851 65962 41860
rect 66168 41064 66220 41070
rect 66168 41006 66220 41012
rect 66180 40905 66208 41006
rect 66166 40896 66222 40905
rect 65654 40828 65962 40837
rect 66166 40831 66222 40840
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40763 65962 40772
rect 65654 39740 65962 39749
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39675 65962 39684
rect 65654 38652 65962 38661
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38587 65962 38596
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 66076 35624 66128 35630
rect 66076 35566 66128 35572
rect 66088 35465 66116 35566
rect 66074 35456 66130 35465
rect 65654 35388 65962 35397
rect 66074 35391 66130 35400
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 67468 33522 67496 44338
rect 67456 33516 67508 33522
rect 67456 33458 67508 33464
rect 65524 33448 65576 33454
rect 65524 33390 65576 33396
rect 66444 33312 66496 33318
rect 66444 33254 66496 33260
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 65800 32972 65852 32978
rect 65800 32914 65852 32920
rect 65812 32434 65840 32914
rect 66168 32836 66220 32842
rect 66168 32778 66220 32784
rect 65984 32768 66036 32774
rect 66180 32745 66208 32778
rect 65984 32710 66036 32716
rect 66166 32736 66222 32745
rect 65996 32502 66024 32710
rect 66166 32671 66222 32680
rect 65984 32496 66036 32502
rect 65984 32438 66036 32444
rect 65800 32428 65852 32434
rect 65800 32370 65852 32376
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 66456 31754 66484 33254
rect 67468 32910 67496 33458
rect 67456 32904 67508 32910
rect 67456 32846 67508 32852
rect 67548 32360 67600 32366
rect 67548 32302 67600 32308
rect 66444 31748 66496 31754
rect 66444 31690 66496 31696
rect 67560 31385 67588 32302
rect 67640 31884 67692 31890
rect 67640 31826 67692 31832
rect 67824 31884 67876 31890
rect 67824 31826 67876 31832
rect 67546 31376 67602 31385
rect 67652 31346 67680 31826
rect 67546 31311 67602 31320
rect 67640 31340 67692 31346
rect 67640 31282 67692 31288
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 66168 30184 66220 30190
rect 66168 30126 66220 30132
rect 66180 30025 66208 30126
rect 66166 30016 66222 30025
rect 65654 29948 65962 29957
rect 66166 29951 66222 29960
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 65524 28484 65576 28490
rect 65524 28426 65576 28432
rect 64788 17128 64840 17134
rect 65536 17105 65564 28426
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 65984 23656 66036 23662
rect 65984 23598 66036 23604
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 64788 17070 64840 17076
rect 65522 17096 65578 17105
rect 63684 11144 63736 11150
rect 63684 11086 63736 11092
rect 59268 8424 59320 8430
rect 59268 8366 59320 8372
rect 56508 3188 56560 3194
rect 56508 3130 56560 3136
rect 59280 1358 59308 8366
rect 64800 4185 64828 17070
rect 65522 17031 65578 17040
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 65996 16574 66024 23598
rect 66168 23248 66220 23254
rect 66166 23216 66168 23225
rect 66220 23216 66222 23225
rect 66166 23151 66222 23160
rect 66076 21480 66128 21486
rect 66076 21422 66128 21428
rect 66088 21185 66116 21422
rect 66074 21176 66130 21185
rect 66074 21111 66130 21120
rect 65996 16546 66116 16574
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 66088 15745 66116 16546
rect 66074 15736 66130 15745
rect 66074 15671 66130 15680
rect 66076 15156 66128 15162
rect 66076 15098 66128 15104
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 66088 14385 66116 15098
rect 66074 14376 66130 14385
rect 66074 14311 66130 14320
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 65248 11688 65300 11694
rect 65248 11630 65300 11636
rect 65260 6225 65288 11630
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 65246 6216 65302 6225
rect 65246 6151 65302 6160
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 64786 4176 64842 4185
rect 64786 4111 64842 4120
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 67836 3534 67864 31826
rect 68928 3596 68980 3602
rect 68928 3538 68980 3544
rect 67824 3528 67876 3534
rect 67824 3470 67876 3476
rect 61200 3460 61252 3466
rect 61200 3402 61252 3408
rect 59268 1352 59320 1358
rect 59268 1294 59320 1300
rect 61212 800 61240 3402
rect 62488 3188 62540 3194
rect 62488 3130 62540 3136
rect 62500 800 62528 3130
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 66168 1352 66220 1358
rect 66168 1294 66220 1300
rect 3422 776 3478 785
rect 3422 711 3478 720
rect 4498 0 4610 800
rect 5786 0 5898 800
rect 7074 0 7186 800
rect 8362 0 8474 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 12226 0 12338 800
rect 13514 0 13626 800
rect 14802 0 14914 800
rect 16090 0 16202 800
rect 17378 0 17490 800
rect 18666 0 18778 800
rect 19954 0 20066 800
rect 21242 0 21354 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 24462 0 24574 800
rect 25750 0 25862 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 29614 0 29726 800
rect 30902 0 31014 800
rect 32190 0 32302 800
rect 33478 0 33590 800
rect 34766 0 34878 800
rect 36054 0 36166 800
rect 37342 0 37454 800
rect 38630 0 38742 800
rect 39918 0 40030 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43782 0 43894 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 47002 0 47114 800
rect 48290 0 48402 800
rect 49578 0 49690 800
rect 50866 0 50978 800
rect 52154 0 52266 800
rect 53442 0 53554 800
rect 54730 0 54842 800
rect 56018 0 56130 800
rect 57306 0 57418 800
rect 58594 0 58706 800
rect 59882 0 59994 800
rect 61170 0 61282 800
rect 62458 0 62570 800
rect 63746 0 63858 800
rect 65034 0 65146 800
rect 66180 785 66208 1294
rect 68940 800 68968 3538
rect 69572 3528 69624 3534
rect 69572 3470 69624 3476
rect 69584 800 69612 3470
rect 66166 776 66222 785
rect 66166 711 66222 720
rect 66322 0 66434 800
rect 67610 0 67722 800
rect 68898 0 69010 800
rect 69542 0 69654 800
<< via2 >>
rect 1490 71440 1546 71496
rect 3514 68720 3570 68776
rect 3422 67360 3478 67416
rect 1398 60596 1400 60616
rect 1400 60596 1452 60616
rect 1452 60596 1454 60616
rect 1398 60560 1454 60596
rect 3330 59200 3386 59256
rect 2778 55120 2834 55176
rect 3330 53760 3386 53816
rect 2962 52400 3018 52456
rect 2870 51040 2926 51096
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4066 49716 4068 49736
rect 4068 49716 4120 49736
rect 4120 49716 4122 49736
rect 4066 49680 4122 49716
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 19580 69658 19636 69660
rect 19660 69658 19716 69660
rect 19740 69658 19796 69660
rect 19820 69658 19876 69660
rect 19580 69606 19626 69658
rect 19626 69606 19636 69658
rect 19660 69606 19690 69658
rect 19690 69606 19702 69658
rect 19702 69606 19716 69658
rect 19740 69606 19754 69658
rect 19754 69606 19766 69658
rect 19766 69606 19796 69658
rect 19820 69606 19830 69658
rect 19830 69606 19876 69658
rect 19580 69604 19636 69606
rect 19660 69604 19716 69606
rect 19740 69604 19796 69606
rect 19820 69604 19876 69606
rect 19580 68570 19636 68572
rect 19660 68570 19716 68572
rect 19740 68570 19796 68572
rect 19820 68570 19876 68572
rect 19580 68518 19626 68570
rect 19626 68518 19636 68570
rect 19660 68518 19690 68570
rect 19690 68518 19702 68570
rect 19702 68518 19716 68570
rect 19740 68518 19754 68570
rect 19754 68518 19766 68570
rect 19766 68518 19796 68570
rect 19820 68518 19830 68570
rect 19830 68518 19876 68570
rect 19580 68516 19636 68518
rect 19660 68516 19716 68518
rect 19740 68516 19796 68518
rect 19820 68516 19876 68518
rect 19580 67482 19636 67484
rect 19660 67482 19716 67484
rect 19740 67482 19796 67484
rect 19820 67482 19876 67484
rect 19580 67430 19626 67482
rect 19626 67430 19636 67482
rect 19660 67430 19690 67482
rect 19690 67430 19702 67482
rect 19702 67430 19716 67482
rect 19740 67430 19754 67482
rect 19754 67430 19766 67482
rect 19766 67430 19796 67482
rect 19820 67430 19830 67482
rect 19830 67430 19876 67482
rect 19580 67428 19636 67430
rect 19660 67428 19716 67430
rect 19740 67428 19796 67430
rect 19820 67428 19876 67430
rect 19580 66394 19636 66396
rect 19660 66394 19716 66396
rect 19740 66394 19796 66396
rect 19820 66394 19876 66396
rect 19580 66342 19626 66394
rect 19626 66342 19636 66394
rect 19660 66342 19690 66394
rect 19690 66342 19702 66394
rect 19702 66342 19716 66394
rect 19740 66342 19754 66394
rect 19754 66342 19766 66394
rect 19766 66342 19796 66394
rect 19820 66342 19830 66394
rect 19830 66342 19876 66394
rect 19580 66340 19636 66342
rect 19660 66340 19716 66342
rect 19740 66340 19796 66342
rect 19820 66340 19876 66342
rect 19580 65306 19636 65308
rect 19660 65306 19716 65308
rect 19740 65306 19796 65308
rect 19820 65306 19876 65308
rect 19580 65254 19626 65306
rect 19626 65254 19636 65306
rect 19660 65254 19690 65306
rect 19690 65254 19702 65306
rect 19702 65254 19716 65306
rect 19740 65254 19754 65306
rect 19754 65254 19766 65306
rect 19766 65254 19796 65306
rect 19820 65254 19830 65306
rect 19830 65254 19876 65306
rect 19580 65252 19636 65254
rect 19660 65252 19716 65254
rect 19740 65252 19796 65254
rect 19820 65252 19876 65254
rect 19580 64218 19636 64220
rect 19660 64218 19716 64220
rect 19740 64218 19796 64220
rect 19820 64218 19876 64220
rect 19580 64166 19626 64218
rect 19626 64166 19636 64218
rect 19660 64166 19690 64218
rect 19690 64166 19702 64218
rect 19702 64166 19716 64218
rect 19740 64166 19754 64218
rect 19754 64166 19766 64218
rect 19766 64166 19796 64218
rect 19820 64166 19830 64218
rect 19830 64166 19876 64218
rect 19580 64164 19636 64166
rect 19660 64164 19716 64166
rect 19740 64164 19796 64166
rect 19820 64164 19876 64166
rect 19580 63130 19636 63132
rect 19660 63130 19716 63132
rect 19740 63130 19796 63132
rect 19820 63130 19876 63132
rect 19580 63078 19626 63130
rect 19626 63078 19636 63130
rect 19660 63078 19690 63130
rect 19690 63078 19702 63130
rect 19702 63078 19716 63130
rect 19740 63078 19754 63130
rect 19754 63078 19766 63130
rect 19766 63078 19796 63130
rect 19820 63078 19830 63130
rect 19830 63078 19876 63130
rect 19580 63076 19636 63078
rect 19660 63076 19716 63078
rect 19740 63076 19796 63078
rect 19820 63076 19876 63078
rect 19580 62042 19636 62044
rect 19660 62042 19716 62044
rect 19740 62042 19796 62044
rect 19820 62042 19876 62044
rect 19580 61990 19626 62042
rect 19626 61990 19636 62042
rect 19660 61990 19690 62042
rect 19690 61990 19702 62042
rect 19702 61990 19716 62042
rect 19740 61990 19754 62042
rect 19754 61990 19766 62042
rect 19766 61990 19796 62042
rect 19820 61990 19830 62042
rect 19830 61990 19876 62042
rect 19580 61988 19636 61990
rect 19660 61988 19716 61990
rect 19740 61988 19796 61990
rect 19820 61988 19876 61990
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4066 47640 4122 47696
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 3054 40840 3110 40896
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 3330 39480 3386 39536
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 3422 38120 3478 38176
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 2870 36760 2926 36816
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 2778 35436 2780 35456
rect 2780 35436 2832 35456
rect 2832 35436 2834 35456
rect 2778 35400 2834 35436
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 3422 31320 3478 31376
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4066 29960 4122 30016
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 3330 22480 3386 22536
rect 3330 15680 3386 15736
rect 3330 12960 3386 13016
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 27276 4068 27296
rect 4068 27276 4120 27296
rect 4120 27276 4122 27296
rect 4066 27240 4122 27276
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4066 25880 4122 25936
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 3974 23840 4030 23896
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 3422 3440 3478 3496
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3606 4800 3662 4856
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3514 2080 3570 2136
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 34940 69114 34996 69116
rect 35020 69114 35076 69116
rect 35100 69114 35156 69116
rect 35180 69114 35236 69116
rect 34940 69062 34986 69114
rect 34986 69062 34996 69114
rect 35020 69062 35050 69114
rect 35050 69062 35062 69114
rect 35062 69062 35076 69114
rect 35100 69062 35114 69114
rect 35114 69062 35126 69114
rect 35126 69062 35156 69114
rect 35180 69062 35190 69114
rect 35190 69062 35236 69114
rect 34940 69060 34996 69062
rect 35020 69060 35076 69062
rect 35100 69060 35156 69062
rect 35180 69060 35236 69062
rect 34940 68026 34996 68028
rect 35020 68026 35076 68028
rect 35100 68026 35156 68028
rect 35180 68026 35236 68028
rect 34940 67974 34986 68026
rect 34986 67974 34996 68026
rect 35020 67974 35050 68026
rect 35050 67974 35062 68026
rect 35062 67974 35076 68026
rect 35100 67974 35114 68026
rect 35114 67974 35126 68026
rect 35126 67974 35156 68026
rect 35180 67974 35190 68026
rect 35190 67974 35236 68026
rect 34940 67972 34996 67974
rect 35020 67972 35076 67974
rect 35100 67972 35156 67974
rect 35180 67972 35236 67974
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 34940 64762 34996 64764
rect 35020 64762 35076 64764
rect 35100 64762 35156 64764
rect 35180 64762 35236 64764
rect 34940 64710 34986 64762
rect 34986 64710 34996 64762
rect 35020 64710 35050 64762
rect 35050 64710 35062 64762
rect 35062 64710 35076 64762
rect 35100 64710 35114 64762
rect 35114 64710 35126 64762
rect 35126 64710 35156 64762
rect 35180 64710 35190 64762
rect 35190 64710 35236 64762
rect 34940 64708 34996 64710
rect 35020 64708 35076 64710
rect 35100 64708 35156 64710
rect 35180 64708 35236 64710
rect 34940 63674 34996 63676
rect 35020 63674 35076 63676
rect 35100 63674 35156 63676
rect 35180 63674 35236 63676
rect 34940 63622 34986 63674
rect 34986 63622 34996 63674
rect 35020 63622 35050 63674
rect 35050 63622 35062 63674
rect 35062 63622 35076 63674
rect 35100 63622 35114 63674
rect 35114 63622 35126 63674
rect 35126 63622 35156 63674
rect 35180 63622 35190 63674
rect 35190 63622 35236 63674
rect 34940 63620 34996 63622
rect 35020 63620 35076 63622
rect 35100 63620 35156 63622
rect 35180 63620 35236 63622
rect 34940 62586 34996 62588
rect 35020 62586 35076 62588
rect 35100 62586 35156 62588
rect 35180 62586 35236 62588
rect 34940 62534 34986 62586
rect 34986 62534 34996 62586
rect 35020 62534 35050 62586
rect 35050 62534 35062 62586
rect 35062 62534 35076 62586
rect 35100 62534 35114 62586
rect 35114 62534 35126 62586
rect 35126 62534 35156 62586
rect 35180 62534 35190 62586
rect 35190 62534 35236 62586
rect 34940 62532 34996 62534
rect 35020 62532 35076 62534
rect 35100 62532 35156 62534
rect 35180 62532 35236 62534
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 69658 50356 69660
rect 50380 69658 50436 69660
rect 50460 69658 50516 69660
rect 50540 69658 50596 69660
rect 50300 69606 50346 69658
rect 50346 69606 50356 69658
rect 50380 69606 50410 69658
rect 50410 69606 50422 69658
rect 50422 69606 50436 69658
rect 50460 69606 50474 69658
rect 50474 69606 50486 69658
rect 50486 69606 50516 69658
rect 50540 69606 50550 69658
rect 50550 69606 50596 69658
rect 50300 69604 50356 69606
rect 50380 69604 50436 69606
rect 50460 69604 50516 69606
rect 50540 69604 50596 69606
rect 50300 68570 50356 68572
rect 50380 68570 50436 68572
rect 50460 68570 50516 68572
rect 50540 68570 50596 68572
rect 50300 68518 50346 68570
rect 50346 68518 50356 68570
rect 50380 68518 50410 68570
rect 50410 68518 50422 68570
rect 50422 68518 50436 68570
rect 50460 68518 50474 68570
rect 50474 68518 50486 68570
rect 50486 68518 50516 68570
rect 50540 68518 50550 68570
rect 50550 68518 50596 68570
rect 50300 68516 50356 68518
rect 50380 68516 50436 68518
rect 50460 68516 50516 68518
rect 50540 68516 50596 68518
rect 50300 67482 50356 67484
rect 50380 67482 50436 67484
rect 50460 67482 50516 67484
rect 50540 67482 50596 67484
rect 50300 67430 50346 67482
rect 50346 67430 50356 67482
rect 50380 67430 50410 67482
rect 50410 67430 50422 67482
rect 50422 67430 50436 67482
rect 50460 67430 50474 67482
rect 50474 67430 50486 67482
rect 50486 67430 50516 67482
rect 50540 67430 50550 67482
rect 50550 67430 50596 67482
rect 50300 67428 50356 67430
rect 50380 67428 50436 67430
rect 50460 67428 50516 67430
rect 50540 67428 50596 67430
rect 50300 66394 50356 66396
rect 50380 66394 50436 66396
rect 50460 66394 50516 66396
rect 50540 66394 50596 66396
rect 50300 66342 50346 66394
rect 50346 66342 50356 66394
rect 50380 66342 50410 66394
rect 50410 66342 50422 66394
rect 50422 66342 50436 66394
rect 50460 66342 50474 66394
rect 50474 66342 50486 66394
rect 50486 66342 50516 66394
rect 50540 66342 50550 66394
rect 50550 66342 50596 66394
rect 50300 66340 50356 66342
rect 50380 66340 50436 66342
rect 50460 66340 50516 66342
rect 50540 66340 50596 66342
rect 50300 65306 50356 65308
rect 50380 65306 50436 65308
rect 50460 65306 50516 65308
rect 50540 65306 50596 65308
rect 50300 65254 50346 65306
rect 50346 65254 50356 65306
rect 50380 65254 50410 65306
rect 50410 65254 50422 65306
rect 50422 65254 50436 65306
rect 50460 65254 50474 65306
rect 50474 65254 50486 65306
rect 50486 65254 50516 65306
rect 50540 65254 50550 65306
rect 50550 65254 50596 65306
rect 50300 65252 50356 65254
rect 50380 65252 50436 65254
rect 50460 65252 50516 65254
rect 50540 65252 50596 65254
rect 50300 64218 50356 64220
rect 50380 64218 50436 64220
rect 50460 64218 50516 64220
rect 50540 64218 50596 64220
rect 50300 64166 50346 64218
rect 50346 64166 50356 64218
rect 50380 64166 50410 64218
rect 50410 64166 50422 64218
rect 50422 64166 50436 64218
rect 50460 64166 50474 64218
rect 50474 64166 50486 64218
rect 50486 64166 50516 64218
rect 50540 64166 50550 64218
rect 50550 64166 50596 64218
rect 50300 64164 50356 64166
rect 50380 64164 50436 64166
rect 50460 64164 50516 64166
rect 50540 64164 50596 64166
rect 50300 63130 50356 63132
rect 50380 63130 50436 63132
rect 50460 63130 50516 63132
rect 50540 63130 50596 63132
rect 50300 63078 50346 63130
rect 50346 63078 50356 63130
rect 50380 63078 50410 63130
rect 50410 63078 50422 63130
rect 50422 63078 50436 63130
rect 50460 63078 50474 63130
rect 50474 63078 50486 63130
rect 50486 63078 50516 63130
rect 50540 63078 50550 63130
rect 50550 63078 50596 63130
rect 50300 63076 50356 63078
rect 50380 63076 50436 63078
rect 50460 63076 50516 63078
rect 50540 63076 50596 63078
rect 50300 62042 50356 62044
rect 50380 62042 50436 62044
rect 50460 62042 50516 62044
rect 50540 62042 50596 62044
rect 50300 61990 50346 62042
rect 50346 61990 50356 62042
rect 50380 61990 50410 62042
rect 50410 61990 50422 62042
rect 50422 61990 50436 62042
rect 50460 61990 50474 62042
rect 50474 61990 50486 62042
rect 50486 61990 50516 62042
rect 50540 61990 50550 62042
rect 50550 61990 50596 62042
rect 50300 61988 50356 61990
rect 50380 61988 50436 61990
rect 50460 61988 50516 61990
rect 50540 61988 50596 61990
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 65660 69114 65716 69116
rect 65740 69114 65796 69116
rect 65820 69114 65876 69116
rect 65900 69114 65956 69116
rect 65660 69062 65706 69114
rect 65706 69062 65716 69114
rect 65740 69062 65770 69114
rect 65770 69062 65782 69114
rect 65782 69062 65796 69114
rect 65820 69062 65834 69114
rect 65834 69062 65846 69114
rect 65846 69062 65876 69114
rect 65900 69062 65910 69114
rect 65910 69062 65956 69114
rect 65660 69060 65716 69062
rect 65740 69060 65796 69062
rect 65820 69060 65876 69062
rect 65900 69060 65956 69062
rect 67454 70080 67510 70136
rect 65660 68026 65716 68028
rect 65740 68026 65796 68028
rect 65820 68026 65876 68028
rect 65900 68026 65956 68028
rect 65660 67974 65706 68026
rect 65706 67974 65716 68026
rect 65740 67974 65770 68026
rect 65770 67974 65782 68026
rect 65782 67974 65796 68026
rect 65820 67974 65834 68026
rect 65834 67974 65846 68026
rect 65846 67974 65876 68026
rect 65900 67974 65910 68026
rect 65910 67974 65956 68026
rect 65660 67972 65716 67974
rect 65740 67972 65796 67974
rect 65820 67972 65876 67974
rect 65900 67972 65956 67974
rect 66166 67360 66222 67416
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 66166 66000 66222 66056
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 65660 64762 65716 64764
rect 65740 64762 65796 64764
rect 65820 64762 65876 64764
rect 65900 64762 65956 64764
rect 65660 64710 65706 64762
rect 65706 64710 65716 64762
rect 65740 64710 65770 64762
rect 65770 64710 65782 64762
rect 65782 64710 65796 64762
rect 65820 64710 65834 64762
rect 65834 64710 65846 64762
rect 65846 64710 65876 64762
rect 65900 64710 65910 64762
rect 65910 64710 65956 64762
rect 65660 64708 65716 64710
rect 65740 64708 65796 64710
rect 65820 64708 65876 64710
rect 65900 64708 65956 64710
rect 65660 63674 65716 63676
rect 65740 63674 65796 63676
rect 65820 63674 65876 63676
rect 65900 63674 65956 63676
rect 65660 63622 65706 63674
rect 65706 63622 65716 63674
rect 65740 63622 65770 63674
rect 65770 63622 65782 63674
rect 65782 63622 65796 63674
rect 65820 63622 65834 63674
rect 65834 63622 65846 63674
rect 65846 63622 65876 63674
rect 65900 63622 65910 63674
rect 65910 63622 65956 63674
rect 65660 63620 65716 63622
rect 65740 63620 65796 63622
rect 65820 63620 65876 63622
rect 65900 63620 65956 63622
rect 65660 62586 65716 62588
rect 65740 62586 65796 62588
rect 65820 62586 65876 62588
rect 65900 62586 65956 62588
rect 65660 62534 65706 62586
rect 65706 62534 65716 62586
rect 65740 62534 65770 62586
rect 65770 62534 65782 62586
rect 65782 62534 65796 62586
rect 65820 62534 65834 62586
rect 65834 62534 65846 62586
rect 65846 62534 65876 62586
rect 65900 62534 65910 62586
rect 65910 62534 65956 62586
rect 65660 62532 65716 62534
rect 65740 62532 65796 62534
rect 65820 62532 65876 62534
rect 65900 62532 65956 62534
rect 66074 61920 66130 61976
rect 65660 61498 65716 61500
rect 65740 61498 65796 61500
rect 65820 61498 65876 61500
rect 65900 61498 65956 61500
rect 65660 61446 65706 61498
rect 65706 61446 65716 61498
rect 65740 61446 65770 61498
rect 65770 61446 65782 61498
rect 65782 61446 65796 61498
rect 65820 61446 65834 61498
rect 65834 61446 65846 61498
rect 65846 61446 65876 61498
rect 65900 61446 65910 61498
rect 65910 61446 65956 61498
rect 65660 61444 65716 61446
rect 65740 61444 65796 61446
rect 65820 61444 65876 61446
rect 65900 61444 65956 61446
rect 66074 60560 66130 60616
rect 65660 60410 65716 60412
rect 65740 60410 65796 60412
rect 65820 60410 65876 60412
rect 65900 60410 65956 60412
rect 65660 60358 65706 60410
rect 65706 60358 65716 60410
rect 65740 60358 65770 60410
rect 65770 60358 65782 60410
rect 65782 60358 65796 60410
rect 65820 60358 65834 60410
rect 65834 60358 65846 60410
rect 65846 60358 65876 60410
rect 65900 60358 65910 60410
rect 65910 60358 65956 60410
rect 65660 60356 65716 60358
rect 65740 60356 65796 60358
rect 65820 60356 65876 60358
rect 65900 60356 65956 60358
rect 64786 59472 64842 59528
rect 66074 59472 66130 59528
rect 64694 56616 64750 56672
rect 65660 59322 65716 59324
rect 65740 59322 65796 59324
rect 65820 59322 65876 59324
rect 65900 59322 65956 59324
rect 65660 59270 65706 59322
rect 65706 59270 65716 59322
rect 65740 59270 65770 59322
rect 65770 59270 65782 59322
rect 65782 59270 65796 59322
rect 65820 59270 65834 59322
rect 65834 59270 65846 59322
rect 65846 59270 65876 59322
rect 65900 59270 65910 59322
rect 65910 59270 65956 59322
rect 65660 59268 65716 59270
rect 65740 59268 65796 59270
rect 65820 59268 65876 59270
rect 65900 59268 65956 59270
rect 65660 58234 65716 58236
rect 65740 58234 65796 58236
rect 65820 58234 65876 58236
rect 65900 58234 65956 58236
rect 65660 58182 65706 58234
rect 65706 58182 65716 58234
rect 65740 58182 65770 58234
rect 65770 58182 65782 58234
rect 65782 58182 65796 58234
rect 65820 58182 65834 58234
rect 65834 58182 65846 58234
rect 65846 58182 65876 58234
rect 65900 58182 65910 58234
rect 65910 58182 65956 58234
rect 65660 58180 65716 58182
rect 65740 58180 65796 58182
rect 65820 58180 65876 58182
rect 65900 58180 65956 58182
rect 66074 57840 66130 57896
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 66074 56616 66130 56672
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 66074 55156 66076 55176
rect 66076 55156 66128 55176
rect 66128 55156 66130 55176
rect 66074 55120 66130 55156
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 67454 63280 67510 63336
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 66074 51040 66130 51096
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 65522 49680 65578 49736
rect 64878 42200 64934 42256
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 67178 46280 67234 46336
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 68098 44940 68154 44976
rect 68098 44920 68100 44940
rect 68100 44920 68152 44940
rect 68152 44920 68154 44940
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 66166 43560 66222 43616
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 66166 40840 66222 40896
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 66074 35400 66130 35456
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 66166 32680 66222 32736
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 67546 31320 67602 31376
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 66166 29960 66222 30016
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 65522 17040 65578 17096
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 66166 23196 66168 23216
rect 66168 23196 66220 23216
rect 66220 23196 66222 23216
rect 66166 23160 66222 23196
rect 66074 21120 66130 21176
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 66074 15680 66130 15736
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 66074 14320 66130 14376
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 65246 6160 65302 6216
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 64786 4120 64842 4176
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 3422 720 3478 776
rect 66166 720 66222 776
<< metal3 >>
rect 0 71498 800 71588
rect 1485 71498 1551 71501
rect 0 71496 1551 71498
rect 0 71440 1490 71496
rect 1546 71440 1551 71496
rect 0 71438 1551 71440
rect 0 71348 800 71438
rect 1485 71435 1551 71438
rect 69200 71348 70000 71588
rect 0 69988 800 70228
rect 67449 70138 67515 70141
rect 69200 70138 70000 70228
rect 67449 70136 70000 70138
rect 67449 70080 67454 70136
rect 67510 70080 70000 70136
rect 67449 70078 70000 70080
rect 67449 70075 67515 70078
rect 69200 69988 70000 70078
rect 19570 69664 19886 69665
rect 19570 69600 19576 69664
rect 19640 69600 19656 69664
rect 19720 69600 19736 69664
rect 19800 69600 19816 69664
rect 19880 69600 19886 69664
rect 19570 69599 19886 69600
rect 50290 69664 50606 69665
rect 50290 69600 50296 69664
rect 50360 69600 50376 69664
rect 50440 69600 50456 69664
rect 50520 69600 50536 69664
rect 50600 69600 50606 69664
rect 50290 69599 50606 69600
rect 4210 69120 4526 69121
rect 4210 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4526 69120
rect 4210 69055 4526 69056
rect 34930 69120 35246 69121
rect 34930 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35246 69120
rect 34930 69055 35246 69056
rect 65650 69120 65966 69121
rect 65650 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65966 69120
rect 65650 69055 65966 69056
rect 0 68778 800 68868
rect 3509 68778 3575 68781
rect 0 68776 3575 68778
rect 0 68720 3514 68776
rect 3570 68720 3575 68776
rect 0 68718 3575 68720
rect 0 68628 800 68718
rect 3509 68715 3575 68718
rect 69200 68628 70000 68868
rect 19570 68576 19886 68577
rect 19570 68512 19576 68576
rect 19640 68512 19656 68576
rect 19720 68512 19736 68576
rect 19800 68512 19816 68576
rect 19880 68512 19886 68576
rect 19570 68511 19886 68512
rect 50290 68576 50606 68577
rect 50290 68512 50296 68576
rect 50360 68512 50376 68576
rect 50440 68512 50456 68576
rect 50520 68512 50536 68576
rect 50600 68512 50606 68576
rect 50290 68511 50606 68512
rect 4210 68032 4526 68033
rect 4210 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4526 68032
rect 4210 67967 4526 67968
rect 34930 68032 35246 68033
rect 34930 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35246 68032
rect 34930 67967 35246 67968
rect 65650 68032 65966 68033
rect 65650 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65966 68032
rect 65650 67967 65966 67968
rect 0 67418 800 67508
rect 19570 67488 19886 67489
rect 19570 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19886 67488
rect 19570 67423 19886 67424
rect 50290 67488 50606 67489
rect 50290 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50606 67488
rect 50290 67423 50606 67424
rect 3417 67418 3483 67421
rect 0 67416 3483 67418
rect 0 67360 3422 67416
rect 3478 67360 3483 67416
rect 0 67358 3483 67360
rect 0 67268 800 67358
rect 3417 67355 3483 67358
rect 66161 67418 66227 67421
rect 69200 67418 70000 67508
rect 66161 67416 70000 67418
rect 66161 67360 66166 67416
rect 66222 67360 70000 67416
rect 66161 67358 70000 67360
rect 66161 67355 66227 67358
rect 69200 67268 70000 67358
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 34930 66944 35246 66945
rect 34930 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35246 66944
rect 34930 66879 35246 66880
rect 65650 66944 65966 66945
rect 65650 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65966 66944
rect 65650 66879 65966 66880
rect 19570 66400 19886 66401
rect 19570 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19886 66400
rect 19570 66335 19886 66336
rect 50290 66400 50606 66401
rect 50290 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50606 66400
rect 50290 66335 50606 66336
rect 0 65908 800 66148
rect 66161 66058 66227 66061
rect 69200 66058 70000 66148
rect 66161 66056 70000 66058
rect 66161 66000 66166 66056
rect 66222 66000 70000 66056
rect 66161 65998 70000 66000
rect 66161 65995 66227 65998
rect 69200 65908 70000 65998
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 34930 65856 35246 65857
rect 34930 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35246 65856
rect 34930 65791 35246 65792
rect 65650 65856 65966 65857
rect 65650 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65966 65856
rect 65650 65791 65966 65792
rect 19570 65312 19886 65313
rect 19570 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19886 65312
rect 19570 65247 19886 65248
rect 50290 65312 50606 65313
rect 50290 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50606 65312
rect 50290 65247 50606 65248
rect 0 64548 800 64788
rect 4210 64768 4526 64769
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 34930 64768 35246 64769
rect 34930 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35246 64768
rect 34930 64703 35246 64704
rect 65650 64768 65966 64769
rect 65650 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65966 64768
rect 65650 64703 65966 64704
rect 69200 64548 70000 64788
rect 19570 64224 19886 64225
rect 19570 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19886 64224
rect 19570 64159 19886 64160
rect 50290 64224 50606 64225
rect 50290 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50606 64224
rect 50290 64159 50606 64160
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 34930 63680 35246 63681
rect 34930 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35246 63680
rect 34930 63615 35246 63616
rect 65650 63680 65966 63681
rect 65650 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65966 63680
rect 65650 63615 65966 63616
rect 0 63188 800 63428
rect 67449 63338 67515 63341
rect 69200 63338 70000 63428
rect 67449 63336 70000 63338
rect 67449 63280 67454 63336
rect 67510 63280 70000 63336
rect 67449 63278 70000 63280
rect 67449 63275 67515 63278
rect 69200 63188 70000 63278
rect 19570 63136 19886 63137
rect 19570 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19886 63136
rect 19570 63071 19886 63072
rect 50290 63136 50606 63137
rect 50290 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50606 63136
rect 50290 63071 50606 63072
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 34930 62592 35246 62593
rect 34930 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35246 62592
rect 34930 62527 35246 62528
rect 65650 62592 65966 62593
rect 65650 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65966 62592
rect 65650 62527 65966 62528
rect 0 61828 800 62068
rect 19570 62048 19886 62049
rect 19570 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19886 62048
rect 19570 61983 19886 61984
rect 50290 62048 50606 62049
rect 50290 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50606 62048
rect 50290 61983 50606 61984
rect 66069 61978 66135 61981
rect 69200 61978 70000 62068
rect 66069 61976 70000 61978
rect 66069 61920 66074 61976
rect 66130 61920 70000 61976
rect 66069 61918 70000 61920
rect 66069 61915 66135 61918
rect 69200 61828 70000 61918
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 34930 61504 35246 61505
rect 34930 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35246 61504
rect 34930 61439 35246 61440
rect 65650 61504 65966 61505
rect 65650 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65966 61504
rect 65650 61439 65966 61440
rect 19570 60960 19886 60961
rect 19570 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19886 60960
rect 19570 60895 19886 60896
rect 50290 60960 50606 60961
rect 50290 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50606 60960
rect 50290 60895 50606 60896
rect 0 60618 800 60708
rect 1393 60618 1459 60621
rect 0 60616 1459 60618
rect 0 60560 1398 60616
rect 1454 60560 1459 60616
rect 0 60558 1459 60560
rect 0 60468 800 60558
rect 1393 60555 1459 60558
rect 66069 60618 66135 60621
rect 69200 60618 70000 60708
rect 66069 60616 70000 60618
rect 66069 60560 66074 60616
rect 66130 60560 70000 60616
rect 66069 60558 70000 60560
rect 66069 60555 66135 60558
rect 69200 60468 70000 60558
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 34930 60416 35246 60417
rect 34930 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35246 60416
rect 34930 60351 35246 60352
rect 65650 60416 65966 60417
rect 65650 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65966 60416
rect 65650 60351 65966 60352
rect 19570 59872 19886 59873
rect 19570 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19886 59872
rect 19570 59807 19886 59808
rect 50290 59872 50606 59873
rect 50290 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50606 59872
rect 50290 59807 50606 59808
rect 64781 59530 64847 59533
rect 66069 59530 66135 59533
rect 64781 59528 66135 59530
rect 64781 59472 64786 59528
rect 64842 59472 66074 59528
rect 66130 59472 66135 59528
rect 64781 59470 66135 59472
rect 64781 59467 64847 59470
rect 66069 59467 66135 59470
rect 0 59258 800 59348
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 34930 59328 35246 59329
rect 34930 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35246 59328
rect 34930 59263 35246 59264
rect 65650 59328 65966 59329
rect 65650 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65966 59328
rect 65650 59263 65966 59264
rect 3325 59258 3391 59261
rect 0 59256 3391 59258
rect 0 59200 3330 59256
rect 3386 59200 3391 59256
rect 0 59198 3391 59200
rect 0 59108 800 59198
rect 3325 59195 3391 59198
rect 69200 59108 70000 59348
rect 19570 58784 19886 58785
rect 19570 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19886 58784
rect 19570 58719 19886 58720
rect 50290 58784 50606 58785
rect 50290 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50606 58784
rect 50290 58719 50606 58720
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 34930 58240 35246 58241
rect 34930 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35246 58240
rect 34930 58175 35246 58176
rect 65650 58240 65966 58241
rect 65650 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65966 58240
rect 65650 58175 65966 58176
rect 0 57748 800 57988
rect 66069 57898 66135 57901
rect 69200 57898 70000 57988
rect 66069 57896 70000 57898
rect 66069 57840 66074 57896
rect 66130 57840 70000 57896
rect 66069 57838 70000 57840
rect 66069 57835 66135 57838
rect 69200 57748 70000 57838
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 65650 57152 65966 57153
rect 65650 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65966 57152
rect 65650 57087 65966 57088
rect 64689 56674 64755 56677
rect 66069 56674 66135 56677
rect 64689 56672 66135 56674
rect 0 56388 800 56628
rect 64689 56616 64694 56672
rect 64750 56616 66074 56672
rect 66130 56616 66135 56672
rect 64689 56614 66135 56616
rect 64689 56611 64755 56614
rect 66069 56611 66135 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 69200 56388 70000 56628
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 65650 56064 65966 56065
rect 65650 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65966 56064
rect 65650 55999 65966 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 0 55178 800 55268
rect 2773 55178 2839 55181
rect 0 55176 2839 55178
rect 0 55120 2778 55176
rect 2834 55120 2839 55176
rect 0 55118 2839 55120
rect 0 55028 800 55118
rect 2773 55115 2839 55118
rect 66069 55178 66135 55181
rect 69200 55178 70000 55268
rect 66069 55176 70000 55178
rect 66069 55120 66074 55176
rect 66130 55120 70000 55176
rect 66069 55118 70000 55120
rect 66069 55115 66135 55118
rect 69200 55028 70000 55118
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 65650 54976 65966 54977
rect 65650 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65966 54976
rect 65650 54911 65966 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 0 53818 800 53908
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 65650 53888 65966 53889
rect 65650 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65966 53888
rect 65650 53823 65966 53824
rect 3325 53818 3391 53821
rect 0 53816 3391 53818
rect 0 53760 3330 53816
rect 3386 53760 3391 53816
rect 0 53758 3391 53760
rect 0 53668 800 53758
rect 3325 53755 3391 53758
rect 69200 53668 70000 53908
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 65650 52800 65966 52801
rect 65650 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65966 52800
rect 65650 52735 65966 52736
rect 0 52458 800 52548
rect 2957 52458 3023 52461
rect 0 52456 3023 52458
rect 0 52400 2962 52456
rect 3018 52400 3023 52456
rect 0 52398 3023 52400
rect 0 52308 800 52398
rect 2957 52395 3023 52398
rect 69200 52308 70000 52548
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 65650 51712 65966 51713
rect 65650 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65966 51712
rect 65650 51647 65966 51648
rect 0 51098 800 51188
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 2865 51098 2931 51101
rect 0 51096 2931 51098
rect 0 51040 2870 51096
rect 2926 51040 2931 51096
rect 0 51038 2931 51040
rect 0 50948 800 51038
rect 2865 51035 2931 51038
rect 66069 51098 66135 51101
rect 69200 51098 70000 51188
rect 66069 51096 70000 51098
rect 66069 51040 66074 51096
rect 66130 51040 70000 51096
rect 66069 51038 70000 51040
rect 66069 51035 66135 51038
rect 69200 50948 70000 51038
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 65650 50624 65966 50625
rect 65650 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65966 50624
rect 65650 50559 65966 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 0 49738 800 49828
rect 4061 49738 4127 49741
rect 0 49736 4127 49738
rect 0 49680 4066 49736
rect 4122 49680 4127 49736
rect 0 49678 4127 49680
rect 0 49588 800 49678
rect 4061 49675 4127 49678
rect 65517 49738 65583 49741
rect 69200 49738 70000 49828
rect 65517 49736 70000 49738
rect 65517 49680 65522 49736
rect 65578 49680 70000 49736
rect 65517 49678 70000 49680
rect 65517 49675 65583 49678
rect 69200 49588 70000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 65650 49536 65966 49537
rect 65650 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65966 49536
rect 65650 49471 65966 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 0 48228 800 48468
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 65650 48448 65966 48449
rect 65650 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65966 48448
rect 65650 48383 65966 48384
rect 69200 48228 70000 48468
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 0 47698 800 47788
rect 4061 47698 4127 47701
rect 0 47696 4127 47698
rect 0 47640 4066 47696
rect 4122 47640 4127 47696
rect 0 47638 4127 47640
rect 0 47548 800 47638
rect 4061 47635 4127 47638
rect 69200 47548 70000 47788
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 65650 47360 65966 47361
rect 65650 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65966 47360
rect 65650 47295 65966 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 0 46188 800 46428
rect 67173 46338 67239 46341
rect 69200 46338 70000 46428
rect 67173 46336 70000 46338
rect 67173 46280 67178 46336
rect 67234 46280 70000 46336
rect 67173 46278 70000 46280
rect 67173 46275 67239 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 65650 46272 65966 46273
rect 65650 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65966 46272
rect 65650 46207 65966 46208
rect 69200 46188 70000 46278
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 65650 45184 65966 45185
rect 65650 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65966 45184
rect 65650 45119 65966 45120
rect 0 44828 800 45068
rect 68093 44978 68159 44981
rect 69200 44978 70000 45068
rect 68093 44976 70000 44978
rect 68093 44920 68098 44976
rect 68154 44920 70000 44976
rect 68093 44918 70000 44920
rect 68093 44915 68159 44918
rect 69200 44828 70000 44918
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 65650 44096 65966 44097
rect 65650 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65966 44096
rect 65650 44031 65966 44032
rect 0 43468 800 43708
rect 66161 43618 66227 43621
rect 69200 43618 70000 43708
rect 66161 43616 70000 43618
rect 66161 43560 66166 43616
rect 66222 43560 70000 43616
rect 66161 43558 70000 43560
rect 66161 43555 66227 43558
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 69200 43468 70000 43558
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 65650 43008 65966 43009
rect 65650 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65966 43008
rect 65650 42943 65966 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 0 42108 800 42348
rect 64873 42258 64939 42261
rect 69200 42258 70000 42348
rect 64873 42256 70000 42258
rect 64873 42200 64878 42256
rect 64934 42200 70000 42256
rect 64873 42198 70000 42200
rect 64873 42195 64939 42198
rect 69200 42108 70000 42198
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 65650 41920 65966 41921
rect 65650 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65966 41920
rect 65650 41855 65966 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 0 40898 800 40988
rect 3049 40898 3115 40901
rect 0 40896 3115 40898
rect 0 40840 3054 40896
rect 3110 40840 3115 40896
rect 0 40838 3115 40840
rect 0 40748 800 40838
rect 3049 40835 3115 40838
rect 66161 40898 66227 40901
rect 69200 40898 70000 40988
rect 66161 40896 70000 40898
rect 66161 40840 66166 40896
rect 66222 40840 70000 40896
rect 66161 40838 70000 40840
rect 66161 40835 66227 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 65650 40832 65966 40833
rect 65650 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65966 40832
rect 65650 40767 65966 40768
rect 69200 40748 70000 40838
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 65650 39744 65966 39745
rect 65650 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65966 39744
rect 65650 39679 65966 39680
rect 0 39538 800 39628
rect 3325 39538 3391 39541
rect 0 39536 3391 39538
rect 0 39480 3330 39536
rect 3386 39480 3391 39536
rect 0 39478 3391 39480
rect 0 39388 800 39478
rect 3325 39475 3391 39478
rect 69200 39388 70000 39628
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 65650 38656 65966 38657
rect 65650 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65966 38656
rect 65650 38591 65966 38592
rect 0 38178 800 38268
rect 3417 38178 3483 38181
rect 0 38176 3483 38178
rect 0 38120 3422 38176
rect 3478 38120 3483 38176
rect 0 38118 3483 38120
rect 0 38028 800 38118
rect 3417 38115 3483 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 69200 38028 70000 38268
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 0 36818 800 36908
rect 2865 36818 2931 36821
rect 0 36816 2931 36818
rect 0 36760 2870 36816
rect 2926 36760 2931 36816
rect 0 36758 2931 36760
rect 0 36668 800 36758
rect 2865 36755 2931 36758
rect 69200 36668 70000 36908
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 0 35458 800 35548
rect 2773 35458 2839 35461
rect 0 35456 2839 35458
rect 0 35400 2778 35456
rect 2834 35400 2839 35456
rect 0 35398 2839 35400
rect 0 35308 800 35398
rect 2773 35395 2839 35398
rect 66069 35458 66135 35461
rect 69200 35458 70000 35548
rect 66069 35456 70000 35458
rect 66069 35400 66074 35456
rect 66130 35400 70000 35456
rect 66069 35398 70000 35400
rect 66069 35395 66135 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 69200 35308 70000 35398
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 0 33948 800 34188
rect 69200 33948 70000 34188
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 0 32588 800 32828
rect 66161 32738 66227 32741
rect 69200 32738 70000 32828
rect 66161 32736 70000 32738
rect 66161 32680 66166 32736
rect 66222 32680 70000 32736
rect 66161 32678 70000 32680
rect 66161 32675 66227 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 69200 32588 70000 32678
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 65650 32063 65966 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 0 31378 800 31468
rect 3417 31378 3483 31381
rect 0 31376 3483 31378
rect 0 31320 3422 31376
rect 3478 31320 3483 31376
rect 0 31318 3483 31320
rect 0 31228 800 31318
rect 3417 31315 3483 31318
rect 67541 31378 67607 31381
rect 69200 31378 70000 31468
rect 67541 31376 70000 31378
rect 67541 31320 67546 31376
rect 67602 31320 70000 31376
rect 67541 31318 70000 31320
rect 67541 31315 67607 31318
rect 69200 31228 70000 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 0 30018 800 30108
rect 4061 30018 4127 30021
rect 0 30016 4127 30018
rect 0 29960 4066 30016
rect 4122 29960 4127 30016
rect 0 29958 4127 29960
rect 0 29868 800 29958
rect 4061 29955 4127 29958
rect 66161 30018 66227 30021
rect 69200 30018 70000 30108
rect 66161 30016 70000 30018
rect 66161 29960 66166 30016
rect 66222 29960 70000 30016
rect 66161 29958 70000 29960
rect 66161 29955 66227 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 69200 29868 70000 29958
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 0 28508 800 28748
rect 69200 28508 70000 28748
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 0 27298 800 27388
rect 4061 27298 4127 27301
rect 0 27296 4127 27298
rect 0 27240 4066 27296
rect 4122 27240 4127 27296
rect 0 27238 4127 27240
rect 0 27148 800 27238
rect 4061 27235 4127 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 69200 27148 70000 27388
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 0 25938 800 26028
rect 4061 25938 4127 25941
rect 0 25936 4127 25938
rect 0 25880 4066 25936
rect 4122 25880 4127 25936
rect 0 25878 4127 25880
rect 0 25788 800 25878
rect 4061 25875 4127 25878
rect 69200 25788 70000 26028
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 0 24428 800 24668
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 69200 24428 70000 24668
rect 0 23898 800 23988
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 3969 23898 4035 23901
rect 0 23896 4035 23898
rect 0 23840 3974 23896
rect 4030 23840 4035 23896
rect 0 23838 4035 23840
rect 0 23748 800 23838
rect 3969 23835 4035 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 66161 23218 66227 23221
rect 69200 23218 70000 23308
rect 66161 23216 70000 23218
rect 66161 23160 66166 23216
rect 66222 23160 70000 23216
rect 66161 23158 70000 23160
rect 66161 23155 66227 23158
rect 69200 23068 70000 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 0 22538 800 22628
rect 3325 22538 3391 22541
rect 0 22536 3391 22538
rect 0 22480 3330 22536
rect 3386 22480 3391 22536
rect 0 22478 3391 22480
rect 0 22388 800 22478
rect 3325 22475 3391 22478
rect 69200 22388 70000 22628
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 0 21028 800 21268
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 66069 21178 66135 21181
rect 69200 21178 70000 21268
rect 66069 21176 70000 21178
rect 66069 21120 66074 21176
rect 66130 21120 70000 21176
rect 66069 21118 70000 21120
rect 66069 21115 66135 21118
rect 69200 21028 70000 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 0 19668 800 19908
rect 69200 19668 70000 19908
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 0 18308 800 18548
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 69200 18308 70000 18548
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 0 16948 800 17188
rect 65517 17098 65583 17101
rect 69200 17098 70000 17188
rect 65517 17096 70000 17098
rect 65517 17040 65522 17096
rect 65578 17040 70000 17096
rect 65517 17038 70000 17040
rect 65517 17035 65583 17038
rect 69200 16948 70000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 0 15738 800 15828
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 3325 15738 3391 15741
rect 0 15736 3391 15738
rect 0 15680 3330 15736
rect 3386 15680 3391 15736
rect 0 15678 3391 15680
rect 0 15588 800 15678
rect 3325 15675 3391 15678
rect 66069 15738 66135 15741
rect 69200 15738 70000 15828
rect 66069 15736 70000 15738
rect 66069 15680 66074 15736
rect 66130 15680 70000 15736
rect 66069 15678 70000 15680
rect 66069 15675 66135 15678
rect 69200 15588 70000 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 0 14228 800 14468
rect 66069 14378 66135 14381
rect 69200 14378 70000 14468
rect 66069 14376 70000 14378
rect 66069 14320 66074 14376
rect 66130 14320 70000 14376
rect 66069 14318 70000 14320
rect 66069 14315 66135 14318
rect 69200 14228 70000 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 0 13018 800 13108
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 3325 13018 3391 13021
rect 0 13016 3391 13018
rect 0 12960 3330 13016
rect 3386 12960 3391 13016
rect 0 12958 3391 12960
rect 0 12868 800 12958
rect 3325 12955 3391 12958
rect 69200 12868 70000 13108
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 0 11508 800 11748
rect 69200 11508 70000 11748
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 0 10148 800 10388
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 69200 10148 70000 10388
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 0 8788 800 9028
rect 69200 8788 70000 9028
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 65650 8127 65966 8128
rect 0 7428 800 7668
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 69200 7428 70000 7668
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 0 6068 800 6308
rect 65241 6218 65307 6221
rect 69200 6218 70000 6308
rect 65241 6216 70000 6218
rect 65241 6160 65246 6216
rect 65302 6160 70000 6216
rect 65241 6158 70000 6160
rect 65241 6155 65307 6158
rect 69200 6068 70000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 0 4858 800 4948
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 3601 4858 3667 4861
rect 69200 4858 70000 4948
rect 0 4856 3667 4858
rect 0 4800 3606 4856
rect 3662 4800 3667 4856
rect 0 4798 3667 4800
rect 0 4708 800 4798
rect 3601 4795 3667 4798
rect 69062 4798 70000 4858
rect 69062 4722 69122 4798
rect 69200 4722 70000 4798
rect 69062 4708 70000 4722
rect 69062 4662 69306 4708
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 64781 4178 64847 4181
rect 69246 4178 69306 4662
rect 64781 4176 69306 4178
rect 64781 4120 64786 4176
rect 64842 4120 69306 4176
rect 64781 4118 69306 4120
rect 64781 4115 64847 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 0 3498 800 3588
rect 3417 3498 3483 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3348 800 3438
rect 3417 3435 3483 3438
rect 69200 3348 70000 3588
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 0 2138 800 2228
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 3509 2138 3575 2141
rect 0 2136 3575 2138
rect 0 2080 3514 2136
rect 3570 2080 3575 2136
rect 0 2078 3575 2080
rect 0 1988 800 2078
rect 3509 2075 3575 2078
rect 69200 1988 70000 2228
rect 0 778 800 868
rect 3417 778 3483 781
rect 0 776 3483 778
rect 0 720 3422 776
rect 3478 720 3483 776
rect 0 718 3483 720
rect 0 628 800 718
rect 3417 715 3483 718
rect 66161 778 66227 781
rect 69200 778 70000 868
rect 66161 776 70000 778
rect 66161 720 66166 776
rect 66222 720 70000 776
rect 66161 718 70000 720
rect 66161 715 66227 718
rect 69200 628 70000 718
<< via3 >>
rect 19576 69660 19640 69664
rect 19576 69604 19580 69660
rect 19580 69604 19636 69660
rect 19636 69604 19640 69660
rect 19576 69600 19640 69604
rect 19656 69660 19720 69664
rect 19656 69604 19660 69660
rect 19660 69604 19716 69660
rect 19716 69604 19720 69660
rect 19656 69600 19720 69604
rect 19736 69660 19800 69664
rect 19736 69604 19740 69660
rect 19740 69604 19796 69660
rect 19796 69604 19800 69660
rect 19736 69600 19800 69604
rect 19816 69660 19880 69664
rect 19816 69604 19820 69660
rect 19820 69604 19876 69660
rect 19876 69604 19880 69660
rect 19816 69600 19880 69604
rect 50296 69660 50360 69664
rect 50296 69604 50300 69660
rect 50300 69604 50356 69660
rect 50356 69604 50360 69660
rect 50296 69600 50360 69604
rect 50376 69660 50440 69664
rect 50376 69604 50380 69660
rect 50380 69604 50436 69660
rect 50436 69604 50440 69660
rect 50376 69600 50440 69604
rect 50456 69660 50520 69664
rect 50456 69604 50460 69660
rect 50460 69604 50516 69660
rect 50516 69604 50520 69660
rect 50456 69600 50520 69604
rect 50536 69660 50600 69664
rect 50536 69604 50540 69660
rect 50540 69604 50596 69660
rect 50596 69604 50600 69660
rect 50536 69600 50600 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 34936 69116 35000 69120
rect 34936 69060 34940 69116
rect 34940 69060 34996 69116
rect 34996 69060 35000 69116
rect 34936 69056 35000 69060
rect 35016 69116 35080 69120
rect 35016 69060 35020 69116
rect 35020 69060 35076 69116
rect 35076 69060 35080 69116
rect 35016 69056 35080 69060
rect 35096 69116 35160 69120
rect 35096 69060 35100 69116
rect 35100 69060 35156 69116
rect 35156 69060 35160 69116
rect 35096 69056 35160 69060
rect 35176 69116 35240 69120
rect 35176 69060 35180 69116
rect 35180 69060 35236 69116
rect 35236 69060 35240 69116
rect 35176 69056 35240 69060
rect 65656 69116 65720 69120
rect 65656 69060 65660 69116
rect 65660 69060 65716 69116
rect 65716 69060 65720 69116
rect 65656 69056 65720 69060
rect 65736 69116 65800 69120
rect 65736 69060 65740 69116
rect 65740 69060 65796 69116
rect 65796 69060 65800 69116
rect 65736 69056 65800 69060
rect 65816 69116 65880 69120
rect 65816 69060 65820 69116
rect 65820 69060 65876 69116
rect 65876 69060 65880 69116
rect 65816 69056 65880 69060
rect 65896 69116 65960 69120
rect 65896 69060 65900 69116
rect 65900 69060 65956 69116
rect 65956 69060 65960 69116
rect 65896 69056 65960 69060
rect 19576 68572 19640 68576
rect 19576 68516 19580 68572
rect 19580 68516 19636 68572
rect 19636 68516 19640 68572
rect 19576 68512 19640 68516
rect 19656 68572 19720 68576
rect 19656 68516 19660 68572
rect 19660 68516 19716 68572
rect 19716 68516 19720 68572
rect 19656 68512 19720 68516
rect 19736 68572 19800 68576
rect 19736 68516 19740 68572
rect 19740 68516 19796 68572
rect 19796 68516 19800 68572
rect 19736 68512 19800 68516
rect 19816 68572 19880 68576
rect 19816 68516 19820 68572
rect 19820 68516 19876 68572
rect 19876 68516 19880 68572
rect 19816 68512 19880 68516
rect 50296 68572 50360 68576
rect 50296 68516 50300 68572
rect 50300 68516 50356 68572
rect 50356 68516 50360 68572
rect 50296 68512 50360 68516
rect 50376 68572 50440 68576
rect 50376 68516 50380 68572
rect 50380 68516 50436 68572
rect 50436 68516 50440 68572
rect 50376 68512 50440 68516
rect 50456 68572 50520 68576
rect 50456 68516 50460 68572
rect 50460 68516 50516 68572
rect 50516 68516 50520 68572
rect 50456 68512 50520 68516
rect 50536 68572 50600 68576
rect 50536 68516 50540 68572
rect 50540 68516 50596 68572
rect 50596 68516 50600 68572
rect 50536 68512 50600 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 34936 68028 35000 68032
rect 34936 67972 34940 68028
rect 34940 67972 34996 68028
rect 34996 67972 35000 68028
rect 34936 67968 35000 67972
rect 35016 68028 35080 68032
rect 35016 67972 35020 68028
rect 35020 67972 35076 68028
rect 35076 67972 35080 68028
rect 35016 67968 35080 67972
rect 35096 68028 35160 68032
rect 35096 67972 35100 68028
rect 35100 67972 35156 68028
rect 35156 67972 35160 68028
rect 35096 67968 35160 67972
rect 35176 68028 35240 68032
rect 35176 67972 35180 68028
rect 35180 67972 35236 68028
rect 35236 67972 35240 68028
rect 35176 67968 35240 67972
rect 65656 68028 65720 68032
rect 65656 67972 65660 68028
rect 65660 67972 65716 68028
rect 65716 67972 65720 68028
rect 65656 67968 65720 67972
rect 65736 68028 65800 68032
rect 65736 67972 65740 68028
rect 65740 67972 65796 68028
rect 65796 67972 65800 68028
rect 65736 67968 65800 67972
rect 65816 68028 65880 68032
rect 65816 67972 65820 68028
rect 65820 67972 65876 68028
rect 65876 67972 65880 68028
rect 65816 67968 65880 67972
rect 65896 68028 65960 68032
rect 65896 67972 65900 68028
rect 65900 67972 65956 68028
rect 65956 67972 65960 68028
rect 65896 67968 65960 67972
rect 19576 67484 19640 67488
rect 19576 67428 19580 67484
rect 19580 67428 19636 67484
rect 19636 67428 19640 67484
rect 19576 67424 19640 67428
rect 19656 67484 19720 67488
rect 19656 67428 19660 67484
rect 19660 67428 19716 67484
rect 19716 67428 19720 67484
rect 19656 67424 19720 67428
rect 19736 67484 19800 67488
rect 19736 67428 19740 67484
rect 19740 67428 19796 67484
rect 19796 67428 19800 67484
rect 19736 67424 19800 67428
rect 19816 67484 19880 67488
rect 19816 67428 19820 67484
rect 19820 67428 19876 67484
rect 19876 67428 19880 67484
rect 19816 67424 19880 67428
rect 50296 67484 50360 67488
rect 50296 67428 50300 67484
rect 50300 67428 50356 67484
rect 50356 67428 50360 67484
rect 50296 67424 50360 67428
rect 50376 67484 50440 67488
rect 50376 67428 50380 67484
rect 50380 67428 50436 67484
rect 50436 67428 50440 67484
rect 50376 67424 50440 67428
rect 50456 67484 50520 67488
rect 50456 67428 50460 67484
rect 50460 67428 50516 67484
rect 50516 67428 50520 67484
rect 50456 67424 50520 67428
rect 50536 67484 50600 67488
rect 50536 67428 50540 67484
rect 50540 67428 50596 67484
rect 50596 67428 50600 67484
rect 50536 67424 50600 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 19576 66396 19640 66400
rect 19576 66340 19580 66396
rect 19580 66340 19636 66396
rect 19636 66340 19640 66396
rect 19576 66336 19640 66340
rect 19656 66396 19720 66400
rect 19656 66340 19660 66396
rect 19660 66340 19716 66396
rect 19716 66340 19720 66396
rect 19656 66336 19720 66340
rect 19736 66396 19800 66400
rect 19736 66340 19740 66396
rect 19740 66340 19796 66396
rect 19796 66340 19800 66396
rect 19736 66336 19800 66340
rect 19816 66396 19880 66400
rect 19816 66340 19820 66396
rect 19820 66340 19876 66396
rect 19876 66340 19880 66396
rect 19816 66336 19880 66340
rect 50296 66396 50360 66400
rect 50296 66340 50300 66396
rect 50300 66340 50356 66396
rect 50356 66340 50360 66396
rect 50296 66336 50360 66340
rect 50376 66396 50440 66400
rect 50376 66340 50380 66396
rect 50380 66340 50436 66396
rect 50436 66340 50440 66396
rect 50376 66336 50440 66340
rect 50456 66396 50520 66400
rect 50456 66340 50460 66396
rect 50460 66340 50516 66396
rect 50516 66340 50520 66396
rect 50456 66336 50520 66340
rect 50536 66396 50600 66400
rect 50536 66340 50540 66396
rect 50540 66340 50596 66396
rect 50596 66340 50600 66396
rect 50536 66336 50600 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 19576 65308 19640 65312
rect 19576 65252 19580 65308
rect 19580 65252 19636 65308
rect 19636 65252 19640 65308
rect 19576 65248 19640 65252
rect 19656 65308 19720 65312
rect 19656 65252 19660 65308
rect 19660 65252 19716 65308
rect 19716 65252 19720 65308
rect 19656 65248 19720 65252
rect 19736 65308 19800 65312
rect 19736 65252 19740 65308
rect 19740 65252 19796 65308
rect 19796 65252 19800 65308
rect 19736 65248 19800 65252
rect 19816 65308 19880 65312
rect 19816 65252 19820 65308
rect 19820 65252 19876 65308
rect 19876 65252 19880 65308
rect 19816 65248 19880 65252
rect 50296 65308 50360 65312
rect 50296 65252 50300 65308
rect 50300 65252 50356 65308
rect 50356 65252 50360 65308
rect 50296 65248 50360 65252
rect 50376 65308 50440 65312
rect 50376 65252 50380 65308
rect 50380 65252 50436 65308
rect 50436 65252 50440 65308
rect 50376 65248 50440 65252
rect 50456 65308 50520 65312
rect 50456 65252 50460 65308
rect 50460 65252 50516 65308
rect 50516 65252 50520 65308
rect 50456 65248 50520 65252
rect 50536 65308 50600 65312
rect 50536 65252 50540 65308
rect 50540 65252 50596 65308
rect 50596 65252 50600 65308
rect 50536 65248 50600 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 34936 64764 35000 64768
rect 34936 64708 34940 64764
rect 34940 64708 34996 64764
rect 34996 64708 35000 64764
rect 34936 64704 35000 64708
rect 35016 64764 35080 64768
rect 35016 64708 35020 64764
rect 35020 64708 35076 64764
rect 35076 64708 35080 64764
rect 35016 64704 35080 64708
rect 35096 64764 35160 64768
rect 35096 64708 35100 64764
rect 35100 64708 35156 64764
rect 35156 64708 35160 64764
rect 35096 64704 35160 64708
rect 35176 64764 35240 64768
rect 35176 64708 35180 64764
rect 35180 64708 35236 64764
rect 35236 64708 35240 64764
rect 35176 64704 35240 64708
rect 65656 64764 65720 64768
rect 65656 64708 65660 64764
rect 65660 64708 65716 64764
rect 65716 64708 65720 64764
rect 65656 64704 65720 64708
rect 65736 64764 65800 64768
rect 65736 64708 65740 64764
rect 65740 64708 65796 64764
rect 65796 64708 65800 64764
rect 65736 64704 65800 64708
rect 65816 64764 65880 64768
rect 65816 64708 65820 64764
rect 65820 64708 65876 64764
rect 65876 64708 65880 64764
rect 65816 64704 65880 64708
rect 65896 64764 65960 64768
rect 65896 64708 65900 64764
rect 65900 64708 65956 64764
rect 65956 64708 65960 64764
rect 65896 64704 65960 64708
rect 19576 64220 19640 64224
rect 19576 64164 19580 64220
rect 19580 64164 19636 64220
rect 19636 64164 19640 64220
rect 19576 64160 19640 64164
rect 19656 64220 19720 64224
rect 19656 64164 19660 64220
rect 19660 64164 19716 64220
rect 19716 64164 19720 64220
rect 19656 64160 19720 64164
rect 19736 64220 19800 64224
rect 19736 64164 19740 64220
rect 19740 64164 19796 64220
rect 19796 64164 19800 64220
rect 19736 64160 19800 64164
rect 19816 64220 19880 64224
rect 19816 64164 19820 64220
rect 19820 64164 19876 64220
rect 19876 64164 19880 64220
rect 19816 64160 19880 64164
rect 50296 64220 50360 64224
rect 50296 64164 50300 64220
rect 50300 64164 50356 64220
rect 50356 64164 50360 64220
rect 50296 64160 50360 64164
rect 50376 64220 50440 64224
rect 50376 64164 50380 64220
rect 50380 64164 50436 64220
rect 50436 64164 50440 64220
rect 50376 64160 50440 64164
rect 50456 64220 50520 64224
rect 50456 64164 50460 64220
rect 50460 64164 50516 64220
rect 50516 64164 50520 64220
rect 50456 64160 50520 64164
rect 50536 64220 50600 64224
rect 50536 64164 50540 64220
rect 50540 64164 50596 64220
rect 50596 64164 50600 64220
rect 50536 64160 50600 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 34936 63676 35000 63680
rect 34936 63620 34940 63676
rect 34940 63620 34996 63676
rect 34996 63620 35000 63676
rect 34936 63616 35000 63620
rect 35016 63676 35080 63680
rect 35016 63620 35020 63676
rect 35020 63620 35076 63676
rect 35076 63620 35080 63676
rect 35016 63616 35080 63620
rect 35096 63676 35160 63680
rect 35096 63620 35100 63676
rect 35100 63620 35156 63676
rect 35156 63620 35160 63676
rect 35096 63616 35160 63620
rect 35176 63676 35240 63680
rect 35176 63620 35180 63676
rect 35180 63620 35236 63676
rect 35236 63620 35240 63676
rect 35176 63616 35240 63620
rect 65656 63676 65720 63680
rect 65656 63620 65660 63676
rect 65660 63620 65716 63676
rect 65716 63620 65720 63676
rect 65656 63616 65720 63620
rect 65736 63676 65800 63680
rect 65736 63620 65740 63676
rect 65740 63620 65796 63676
rect 65796 63620 65800 63676
rect 65736 63616 65800 63620
rect 65816 63676 65880 63680
rect 65816 63620 65820 63676
rect 65820 63620 65876 63676
rect 65876 63620 65880 63676
rect 65816 63616 65880 63620
rect 65896 63676 65960 63680
rect 65896 63620 65900 63676
rect 65900 63620 65956 63676
rect 65956 63620 65960 63676
rect 65896 63616 65960 63620
rect 19576 63132 19640 63136
rect 19576 63076 19580 63132
rect 19580 63076 19636 63132
rect 19636 63076 19640 63132
rect 19576 63072 19640 63076
rect 19656 63132 19720 63136
rect 19656 63076 19660 63132
rect 19660 63076 19716 63132
rect 19716 63076 19720 63132
rect 19656 63072 19720 63076
rect 19736 63132 19800 63136
rect 19736 63076 19740 63132
rect 19740 63076 19796 63132
rect 19796 63076 19800 63132
rect 19736 63072 19800 63076
rect 19816 63132 19880 63136
rect 19816 63076 19820 63132
rect 19820 63076 19876 63132
rect 19876 63076 19880 63132
rect 19816 63072 19880 63076
rect 50296 63132 50360 63136
rect 50296 63076 50300 63132
rect 50300 63076 50356 63132
rect 50356 63076 50360 63132
rect 50296 63072 50360 63076
rect 50376 63132 50440 63136
rect 50376 63076 50380 63132
rect 50380 63076 50436 63132
rect 50436 63076 50440 63132
rect 50376 63072 50440 63076
rect 50456 63132 50520 63136
rect 50456 63076 50460 63132
rect 50460 63076 50516 63132
rect 50516 63076 50520 63132
rect 50456 63072 50520 63076
rect 50536 63132 50600 63136
rect 50536 63076 50540 63132
rect 50540 63076 50596 63132
rect 50596 63076 50600 63132
rect 50536 63072 50600 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 34936 62588 35000 62592
rect 34936 62532 34940 62588
rect 34940 62532 34996 62588
rect 34996 62532 35000 62588
rect 34936 62528 35000 62532
rect 35016 62588 35080 62592
rect 35016 62532 35020 62588
rect 35020 62532 35076 62588
rect 35076 62532 35080 62588
rect 35016 62528 35080 62532
rect 35096 62588 35160 62592
rect 35096 62532 35100 62588
rect 35100 62532 35156 62588
rect 35156 62532 35160 62588
rect 35096 62528 35160 62532
rect 35176 62588 35240 62592
rect 35176 62532 35180 62588
rect 35180 62532 35236 62588
rect 35236 62532 35240 62588
rect 35176 62528 35240 62532
rect 65656 62588 65720 62592
rect 65656 62532 65660 62588
rect 65660 62532 65716 62588
rect 65716 62532 65720 62588
rect 65656 62528 65720 62532
rect 65736 62588 65800 62592
rect 65736 62532 65740 62588
rect 65740 62532 65796 62588
rect 65796 62532 65800 62588
rect 65736 62528 65800 62532
rect 65816 62588 65880 62592
rect 65816 62532 65820 62588
rect 65820 62532 65876 62588
rect 65876 62532 65880 62588
rect 65816 62528 65880 62532
rect 65896 62588 65960 62592
rect 65896 62532 65900 62588
rect 65900 62532 65956 62588
rect 65956 62532 65960 62588
rect 65896 62528 65960 62532
rect 19576 62044 19640 62048
rect 19576 61988 19580 62044
rect 19580 61988 19636 62044
rect 19636 61988 19640 62044
rect 19576 61984 19640 61988
rect 19656 62044 19720 62048
rect 19656 61988 19660 62044
rect 19660 61988 19716 62044
rect 19716 61988 19720 62044
rect 19656 61984 19720 61988
rect 19736 62044 19800 62048
rect 19736 61988 19740 62044
rect 19740 61988 19796 62044
rect 19796 61988 19800 62044
rect 19736 61984 19800 61988
rect 19816 62044 19880 62048
rect 19816 61988 19820 62044
rect 19820 61988 19876 62044
rect 19876 61988 19880 62044
rect 19816 61984 19880 61988
rect 50296 62044 50360 62048
rect 50296 61988 50300 62044
rect 50300 61988 50356 62044
rect 50356 61988 50360 62044
rect 50296 61984 50360 61988
rect 50376 62044 50440 62048
rect 50376 61988 50380 62044
rect 50380 61988 50436 62044
rect 50436 61988 50440 62044
rect 50376 61984 50440 61988
rect 50456 62044 50520 62048
rect 50456 61988 50460 62044
rect 50460 61988 50516 62044
rect 50516 61988 50520 62044
rect 50456 61984 50520 61988
rect 50536 62044 50600 62048
rect 50536 61988 50540 62044
rect 50540 61988 50596 62044
rect 50596 61988 50600 62044
rect 50536 61984 50600 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 65656 61500 65720 61504
rect 65656 61444 65660 61500
rect 65660 61444 65716 61500
rect 65716 61444 65720 61500
rect 65656 61440 65720 61444
rect 65736 61500 65800 61504
rect 65736 61444 65740 61500
rect 65740 61444 65796 61500
rect 65796 61444 65800 61500
rect 65736 61440 65800 61444
rect 65816 61500 65880 61504
rect 65816 61444 65820 61500
rect 65820 61444 65876 61500
rect 65876 61444 65880 61500
rect 65816 61440 65880 61444
rect 65896 61500 65960 61504
rect 65896 61444 65900 61500
rect 65900 61444 65956 61500
rect 65956 61444 65960 61500
rect 65896 61440 65960 61444
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 65656 60412 65720 60416
rect 65656 60356 65660 60412
rect 65660 60356 65716 60412
rect 65716 60356 65720 60412
rect 65656 60352 65720 60356
rect 65736 60412 65800 60416
rect 65736 60356 65740 60412
rect 65740 60356 65796 60412
rect 65796 60356 65800 60412
rect 65736 60352 65800 60356
rect 65816 60412 65880 60416
rect 65816 60356 65820 60412
rect 65820 60356 65876 60412
rect 65876 60356 65880 60412
rect 65816 60352 65880 60356
rect 65896 60412 65960 60416
rect 65896 60356 65900 60412
rect 65900 60356 65956 60412
rect 65956 60356 65960 60412
rect 65896 60352 65960 60356
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 65656 59324 65720 59328
rect 65656 59268 65660 59324
rect 65660 59268 65716 59324
rect 65716 59268 65720 59324
rect 65656 59264 65720 59268
rect 65736 59324 65800 59328
rect 65736 59268 65740 59324
rect 65740 59268 65796 59324
rect 65796 59268 65800 59324
rect 65736 59264 65800 59268
rect 65816 59324 65880 59328
rect 65816 59268 65820 59324
rect 65820 59268 65876 59324
rect 65876 59268 65880 59324
rect 65816 59264 65880 59268
rect 65896 59324 65960 59328
rect 65896 59268 65900 59324
rect 65900 59268 65956 59324
rect 65956 59268 65960 59324
rect 65896 59264 65960 59268
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 65656 58236 65720 58240
rect 65656 58180 65660 58236
rect 65660 58180 65716 58236
rect 65716 58180 65720 58236
rect 65656 58176 65720 58180
rect 65736 58236 65800 58240
rect 65736 58180 65740 58236
rect 65740 58180 65796 58236
rect 65796 58180 65800 58236
rect 65736 58176 65800 58180
rect 65816 58236 65880 58240
rect 65816 58180 65820 58236
rect 65820 58180 65876 58236
rect 65876 58180 65880 58236
rect 65816 58176 65880 58180
rect 65896 58236 65960 58240
rect 65896 58180 65900 58236
rect 65900 58180 65956 58236
rect 65956 58180 65960 58236
rect 65896 58176 65960 58180
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 69120 4528 69680
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 65856 4528 66880
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 69664 19888 69680
rect 19568 69600 19576 69664
rect 19640 69600 19656 69664
rect 19720 69600 19736 69664
rect 19800 69600 19816 69664
rect 19880 69600 19888 69664
rect 19568 68576 19888 69600
rect 19568 68512 19576 68576
rect 19640 68512 19656 68576
rect 19720 68512 19736 68576
rect 19800 68512 19816 68576
rect 19880 68512 19888 68576
rect 19568 67488 19888 68512
rect 19568 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19888 67488
rect 19568 66400 19888 67424
rect 19568 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19888 66400
rect 19568 65312 19888 66336
rect 19568 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19888 65312
rect 19568 64224 19888 65248
rect 19568 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19888 64224
rect 19568 63136 19888 64160
rect 19568 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19888 63136
rect 19568 62048 19888 63072
rect 19568 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19888 62048
rect 19568 60960 19888 61984
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 59872 19888 60896
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 69120 35248 69680
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 68032 35248 69056
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 66944 35248 67968
rect 34928 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35248 66944
rect 34928 65856 35248 66880
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 64768 35248 65792
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 63680 35248 64704
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 62592 35248 63616
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 61504 35248 62528
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59328 35248 60352
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 69664 50608 69680
rect 50288 69600 50296 69664
rect 50360 69600 50376 69664
rect 50440 69600 50456 69664
rect 50520 69600 50536 69664
rect 50600 69600 50608 69664
rect 50288 68576 50608 69600
rect 50288 68512 50296 68576
rect 50360 68512 50376 68576
rect 50440 68512 50456 68576
rect 50520 68512 50536 68576
rect 50600 68512 50608 68576
rect 50288 67488 50608 68512
rect 50288 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50608 67488
rect 50288 66400 50608 67424
rect 50288 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50608 66400
rect 50288 65312 50608 66336
rect 50288 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50608 65312
rect 50288 64224 50608 65248
rect 50288 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50608 64224
rect 50288 63136 50608 64160
rect 50288 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50608 63136
rect 50288 62048 50608 63072
rect 50288 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50608 62048
rect 50288 60960 50608 61984
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 69120 65968 69680
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 68032 65968 69056
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 66944 65968 67968
rect 65648 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65968 66944
rect 65648 65856 65968 66880
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 64768 65968 65792
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 63680 65968 64704
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 62592 65968 63616
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 61504 65968 62528
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 60416 65968 61440
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 59328 65968 60352
rect 65648 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65968 59328
rect 65648 58240 65968 59264
rect 65648 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65968 58240
rect 65648 57152 65968 58176
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 30636 0 1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1649977179
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_285 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_292
timestamp 1649977179
transform 1 0 27968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1649977179
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1649977179
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1649977179
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1649977179
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1649977179
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1649977179
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1649977179
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1649977179
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_424 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1649977179
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1649977179
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1649977179
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1649977179
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1649977179
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1649977179
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1649977179
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1649977179
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1649977179
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1649977179
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1649977179
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1649977179
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1649977179
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1649977179
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1649977179
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1649977179
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1649977179
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1649977179
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1649977179
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1649977179
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1649977179
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1649977179
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1649977179
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1649977179
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1649977179
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1649977179
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1649977179
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1649977179
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1649977179
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729
timestamp 1649977179
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1649977179
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_284
timestamp 1649977179
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_309
timestamp 1649977179
transform 1 0 29532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_321
timestamp 1649977179
transform 1 0 30636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1649977179
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1649977179
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1649977179
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_412
timestamp 1649977179
transform 1 0 39008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_437
timestamp 1649977179
transform 1 0 41308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1649977179
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1649977179
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1649977179
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1649977179
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1649977179
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1649977179
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1649977179
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1649977179
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1649977179
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1649977179
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1649977179
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1649977179
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1649977179
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1649977179
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1649977179
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1649977179
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1649977179
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1649977179
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1649977179
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1649977179
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1649977179
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1649977179
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1649977179
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1649977179
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1649977179
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1649977179
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1649977179
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1649977179
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1649977179
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1649977179
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_421 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_429
timestamp 1649977179
transform 1 0 40572 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_451
timestamp 1649977179
transform 1 0 42596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_463
timestamp 1649977179
transform 1 0 43700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1649977179
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1649977179
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1649977179
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1649977179
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1649977179
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1649977179
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1649977179
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1649977179
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1649977179
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1649977179
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1649977179
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1649977179
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1649977179
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1649977179
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1649977179
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1649977179
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1649977179
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1649977179
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1649977179
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1649977179
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1649977179
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1649977179
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_725
timestamp 1649977179
transform 1 0 67804 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1649977179
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1649977179
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1649977179
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1649977179
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1649977179
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1649977179
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1649977179
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1649977179
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1649977179
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1649977179
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1649977179
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_729
timestamp 1649977179
transform 1 0 68172 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1649977179
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1649977179
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1649977179
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1649977179
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1649977179
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1649977179
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1649977179
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1649977179
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1649977179
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1649977179
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1649977179
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1649977179
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1649977179
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_725
timestamp 1649977179
transform 1 0 67804 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1649977179
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1649977179
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1649977179
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1649977179
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1649977179
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1649977179
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1649977179
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1649977179
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1649977179
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1649977179
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1649977179
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1649977179
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1649977179
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1649977179
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1649977179
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_729
timestamp 1649977179
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1649977179
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1649977179
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1649977179
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1649977179
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1649977179
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1649977179
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1649977179
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1649977179
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1649977179
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1649977179
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1649977179
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_725
timestamp 1649977179
transform 1 0 67804 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1649977179
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1649977179
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1649977179
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1649977179
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1649977179
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1649977179
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1649977179
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1649977179
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1649977179
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1649977179
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1649977179
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_729
timestamp 1649977179
transform 1 0 68172 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1649977179
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1649977179
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1649977179
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1649977179
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1649977179
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1649977179
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1649977179
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1649977179
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1649977179
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1649977179
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1649977179
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_725
timestamp 1649977179
transform 1 0 67804 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1649977179
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1649977179
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1649977179
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1649977179
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1649977179
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1649977179
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1649977179
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1649977179
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1649977179
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1649977179
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1649977179
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1649977179
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_729
timestamp 1649977179
transform 1 0 68172 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1649977179
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1649977179
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1649977179
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1649977179
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1649977179
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1649977179
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1649977179
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1649977179
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1649977179
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1649977179
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1649977179
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_725
timestamp 1649977179
transform 1 0 67804 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_284
timestamp 1649977179
transform 1 0 27232 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_296
timestamp 1649977179
transform 1 0 28336 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_308
timestamp 1649977179
transform 1 0 29440 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_320
timestamp 1649977179
transform 1 0 30544 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1649977179
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_581 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 54556 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_604
timestamp 1649977179
transform 1 0 56672 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1649977179
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1649977179
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1649977179
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1649977179
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1649977179
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1649977179
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1649977179
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1649977179
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1649977179
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1649977179
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1649977179
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_729
timestamp 1649977179
transform 1 0 68172 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1649977179
transform 1 0 26036 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_296
timestamp 1649977179
transform 1 0 28336 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_462
timestamp 1649977179
transform 1 0 43608 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_474
timestamp 1649977179
transform 1 0 44712 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_577
timestamp 1649977179
transform 1 0 54188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_582
timestamp 1649977179
transform 1 0 54648 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_592
timestamp 1649977179
transform 1 0 55568 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_604
timestamp 1649977179
transform 1 0 56672 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_616
timestamp 1649977179
transform 1 0 57776 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_628
timestamp 1649977179
transform 1 0 58880 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_640
timestamp 1649977179
transform 1 0 59984 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1649977179
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1649977179
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1649977179
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1649977179
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1649977179
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1649977179
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1649977179
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1649977179
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_725
timestamp 1649977179
transform 1 0 67804 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1649977179
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_457
timestamp 1649977179
transform 1 0 43148 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_479
timestamp 1649977179
transform 1 0 45172 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_491
timestamp 1649977179
transform 1 0 46276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1649977179
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1649977179
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1649977179
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1649977179
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1649977179
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1649977179
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1649977179
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1649977179
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1649977179
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1649977179
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1649977179
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_729
timestamp 1649977179
transform 1 0 68172 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_292
timestamp 1649977179
transform 1 0 27968 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1649977179
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1649977179
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_462
timestamp 1649977179
transform 1 0 43608 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_474
timestamp 1649977179
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1649977179
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1649977179
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1649977179
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1649977179
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1649977179
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1649977179
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1649977179
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1649977179
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1649977179
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1649977179
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1649977179
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_725
timestamp 1649977179
transform 1 0 67804 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_257
timestamp 1649977179
transform 1 0 24748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_263
timestamp 1649977179
transform 1 0 25300 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_271
timestamp 1649977179
transform 1 0 26036 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1649977179
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_323
timestamp 1649977179
transform 1 0 30820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_369
timestamp 1649977179
transform 1 0 35052 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1649977179
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1649977179
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1649977179
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1649977179
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1649977179
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1649977179
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1649977179
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1649977179
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1649977179
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1649977179
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1649977179
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_729
timestamp 1649977179
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_276
timestamp 1649977179
transform 1 0 26496 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_283
timestamp 1649977179
transform 1 0 27140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_295
timestamp 1649977179
transform 1 0 28244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_336
timestamp 1649977179
transform 1 0 32016 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_348
timestamp 1649977179
transform 1 0 33120 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_356
timestamp 1649977179
transform 1 0 33856 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1649977179
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_388
timestamp 1649977179
transform 1 0 36800 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_400
timestamp 1649977179
transform 1 0 37904 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_412
timestamp 1649977179
transform 1 0 39008 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1649977179
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1649977179
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1649977179
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1649977179
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1649977179
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_669
timestamp 1649977179
transform 1 0 62652 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_678
timestamp 1649977179
transform 1 0 63480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_690
timestamp 1649977179
transform 1 0 64584 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_698
timestamp 1649977179
transform 1 0 65320 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1649977179
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1649977179
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_725
timestamp 1649977179
transform 1 0 67804 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_258
timestamp 1649977179
transform 1 0 24840 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_270
timestamp 1649977179
transform 1 0 25944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1649977179
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_313
timestamp 1649977179
transform 1 0 29900 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_318
timestamp 1649977179
transform 1 0 30360 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_330
timestamp 1649977179
transform 1 0 31464 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_356
timestamp 1649977179
transform 1 0 33856 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_381
timestamp 1649977179
transform 1 0 36156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_389
timestamp 1649977179
transform 1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1649977179
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1649977179
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1649977179
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1649977179
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1649977179
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1649977179
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1649977179
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1649977179
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_673
timestamp 1649977179
transform 1 0 63020 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_698
timestamp 1649977179
transform 1 0 65320 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_710
timestamp 1649977179
transform 1 0 66424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_722
timestamp 1649977179
transform 1 0 67528 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_729
timestamp 1649977179
transform 1 0 68172 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_368
timestamp 1649977179
transform 1 0 34960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_372
timestamp 1649977179
transform 1 0 35328 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_394
timestamp 1649977179
transform 1 0 37352 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_406
timestamp 1649977179
transform 1 0 38456 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_418
timestamp 1649977179
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1649977179
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1649977179
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1649977179
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1649977179
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1649977179
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_669
timestamp 1649977179
transform 1 0 62652 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_680
timestamp 1649977179
transform 1 0 63664 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_692
timestamp 1649977179
transform 1 0 64768 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1649977179
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1649977179
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_725
timestamp 1649977179
transform 1 0 67804 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_377
timestamp 1649977179
transform 1 0 35788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1649977179
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1649977179
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1649977179
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1649977179
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1649977179
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1649977179
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1649977179
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1649977179
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1649977179
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1649977179
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1649977179
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1649977179
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_729
timestamp 1649977179
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1649977179
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_207
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_219
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_230
timestamp 1649977179
transform 1 0 22264 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_242
timestamp 1649977179
transform 1 0 23368 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1649977179
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_373
timestamp 1649977179
transform 1 0 35420 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1649977179
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1649977179
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1649977179
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1649977179
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1649977179
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1649977179
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1649977179
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1649977179
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1649977179
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1649977179
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1649977179
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_725
timestamp 1649977179
transform 1 0 67804 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1649977179
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_248
timestamp 1649977179
transform 1 0 23920 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_260
timestamp 1649977179
transform 1 0 25024 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_272
timestamp 1649977179
transform 1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1649977179
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1649977179
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1649977179
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1649977179
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1649977179
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1649977179
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1649977179
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1649977179
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1649977179
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1649977179
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1649977179
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_729
timestamp 1649977179
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_130
timestamp 1649977179
transform 1 0 13064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_202
timestamp 1649977179
transform 1 0 19688 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_214
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_226
timestamp 1649977179
transform 1 0 21896 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_231
timestamp 1649977179
transform 1 0 22356 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1649977179
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1649977179
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1649977179
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1649977179
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1649977179
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1649977179
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1649977179
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1649977179
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1649977179
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1649977179
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1649977179
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1649977179
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_725
timestamp 1649977179
transform 1 0 67804 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_148
timestamp 1649977179
transform 1 0 14720 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_160
timestamp 1649977179
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1649977179
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1649977179
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1649977179
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1649977179
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1649977179
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1649977179
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1649977179
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1649977179
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1649977179
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1649977179
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1649977179
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_729
timestamp 1649977179
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_127
timestamp 1649977179
transform 1 0 12788 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_131
timestamp 1649977179
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1649977179
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1649977179
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1649977179
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1649977179
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1649977179
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1649977179
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1649977179
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1649977179
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1649977179
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1649977179
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1649977179
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_725
timestamp 1649977179
transform 1 0 67804 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1649977179
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1649977179
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1649977179
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1649977179
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1649977179
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1649977179
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1649977179
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1649977179
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1649977179
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1649977179
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1649977179
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_729
timestamp 1649977179
transform 1 0 68172 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1649977179
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1649977179
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1649977179
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1649977179
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1649977179
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1649977179
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1649977179
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1649977179
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1649977179
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1649977179
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1649977179
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_725
timestamp 1649977179
transform 1 0 67804 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1649977179
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1649977179
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1649977179
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1649977179
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1649977179
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1649977179
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1649977179
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1649977179
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1649977179
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_694
timestamp 1649977179
transform 1 0 64952 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_706
timestamp 1649977179
transform 1 0 66056 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_718
timestamp 1649977179
transform 1 0 67160 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_726
timestamp 1649977179
transform 1 0 67896 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_729
timestamp 1649977179
transform 1 0 68172 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1649977179
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1649977179
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1649977179
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1649977179
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1649977179
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1649977179
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_672
timestamp 1649977179
transform 1 0 62928 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_679
timestamp 1649977179
transform 1 0 63572 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_691
timestamp 1649977179
transform 1 0 64676 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1649977179
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1649977179
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1649977179
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_725
timestamp 1649977179
transform 1 0 67804 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_48
timestamp 1649977179
transform 1 0 5520 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1649977179
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1649977179
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1649977179
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1649977179
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1649977179
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1649977179
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1649977179
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1649977179
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1649977179
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1649977179
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1649977179
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1649977179
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_729
timestamp 1649977179
transform 1 0 68172 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_339
timestamp 1649977179
transform 1 0 32292 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_343
timestamp 1649977179
transform 1 0 32660 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_355
timestamp 1649977179
transform 1 0 33764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1649977179
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1649977179
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1649977179
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1649977179
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1649977179
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1649977179
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1649977179
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1649977179
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1649977179
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1649977179
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1649977179
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1649977179
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1649977179
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1649977179
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1649977179
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_725
timestamp 1649977179
transform 1 0 67804 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_358
timestamp 1649977179
transform 1 0 34040 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_370
timestamp 1649977179
transform 1 0 35144 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_382
timestamp 1649977179
transform 1 0 36248 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1649977179
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1649977179
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1649977179
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1649977179
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1649977179
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1649977179
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1649977179
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1649977179
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1649977179
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1649977179
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1649977179
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1649977179
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1649977179
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1649977179
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_729
timestamp 1649977179
transform 1 0 68172 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_340
timestamp 1649977179
transform 1 0 32384 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_352
timestamp 1649977179
transform 1 0 33488 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1649977179
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1649977179
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1649977179
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1649977179
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1649977179
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1649977179
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1649977179
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1649977179
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1649977179
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1649977179
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1649977179
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_725
timestamp 1649977179
transform 1 0 67804 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1649977179
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1649977179
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1649977179
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1649977179
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1649977179
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1649977179
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1649977179
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1649977179
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1649977179
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1649977179
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1649977179
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_729
timestamp 1649977179
transform 1 0 68172 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1649977179
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1649977179
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1649977179
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1649977179
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1649977179
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_669
timestamp 1649977179
transform 1 0 62652 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_673
timestamp 1649977179
transform 1 0 63020 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_677
timestamp 1649977179
transform 1 0 63388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_689
timestamp 1649977179
transform 1 0 64492 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_697
timestamp 1649977179
transform 1 0 65228 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1649977179
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1649977179
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_725
timestamp 1649977179
transform 1 0 67804 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1649977179
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1649977179
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1649977179
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1649977179
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1649977179
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1649977179
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1649977179
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1649977179
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_673
timestamp 1649977179
transform 1 0 63020 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_695
timestamp 1649977179
transform 1 0 65044 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_707
timestamp 1649977179
transform 1 0 66148 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_719
timestamp 1649977179
transform 1 0 67252 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1649977179
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_729
timestamp 1649977179
transform 1 0 68172 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_58
timestamp 1649977179
transform 1 0 6440 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_70
timestamp 1649977179
transform 1 0 7544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1649977179
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_124
timestamp 1649977179
transform 1 0 12512 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1649977179
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1649977179
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_556
timestamp 1649977179
transform 1 0 52256 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_568
timestamp 1649977179
transform 1 0 53360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_580
timestamp 1649977179
transform 1 0 54464 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1649977179
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1649977179
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1649977179
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1649977179
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1649977179
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_669
timestamp 1649977179
transform 1 0 62652 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_675
timestamp 1649977179
transform 1 0 63204 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_687
timestamp 1649977179
transform 1 0 64308 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1649977179
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1649977179
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1649977179
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_725
timestamp 1649977179
transform 1 0 67804 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_35
timestamp 1649977179
transform 1 0 4324 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_40
timestamp 1649977179
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1649977179
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1649977179
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1649977179
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_540
timestamp 1649977179
transform 1 0 50784 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_547
timestamp 1649977179
transform 1 0 51428 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1649977179
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_641
timestamp 1649977179
transform 1 0 60076 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_668
timestamp 1649977179
transform 1 0 62560 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1649977179
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1649977179
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1649977179
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1649977179
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1649977179
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1649977179
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_729
timestamp 1649977179
transform 1 0 68172 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_108
timestamp 1649977179
transform 1 0 11040 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_115
timestamp 1649977179
transform 1 0 11684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_127
timestamp 1649977179
transform 1 0 12788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_620
timestamp 1649977179
transform 1 0 58144 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_632
timestamp 1649977179
transform 1 0 59248 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_645
timestamp 1649977179
transform 1 0 60444 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_651
timestamp 1649977179
transform 1 0 60996 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_658
timestamp 1649977179
transform 1 0 61640 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_670
timestamp 1649977179
transform 1 0 62744 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_682
timestamp 1649977179
transform 1 0 63848 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_694
timestamp 1649977179
transform 1 0 64952 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1649977179
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1649977179
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_725
timestamp 1649977179
transform 1 0 67804 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1649977179
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1649977179
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1649977179
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1649977179
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1649977179
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1649977179
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1649977179
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1649977179
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1649977179
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1649977179
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_729
timestamp 1649977179
transform 1 0 68172 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_624
timestamp 1649977179
transform 1 0 58512 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_636
timestamp 1649977179
transform 1 0 59616 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1649977179
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1649977179
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1649977179
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1649977179
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1649977179
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1649977179
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1649977179
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1649977179
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_725
timestamp 1649977179
transform 1 0 67804 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_297
timestamp 1649977179
transform 1 0 28428 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_304
timestamp 1649977179
transform 1 0 29072 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_316
timestamp 1649977179
transform 1 0 30176 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_328
timestamp 1649977179
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_367
timestamp 1649977179
transform 1 0 34868 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_371
timestamp 1649977179
transform 1 0 35236 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_383
timestamp 1649977179
transform 1 0 36340 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1649977179
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1649977179
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1649977179
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1649977179
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1649977179
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1649977179
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1649977179
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1649977179
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1649977179
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1649977179
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1649977179
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1649977179
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_729
timestamp 1649977179
transform 1 0 68172 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_388
timestamp 1649977179
transform 1 0 36800 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_400
timestamp 1649977179
transform 1 0 37904 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_412
timestamp 1649977179
transform 1 0 39008 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1649977179
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1649977179
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1649977179
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1649977179
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1649977179
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1649977179
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1649977179
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1649977179
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1649977179
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1649977179
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1649977179
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_725
timestamp 1649977179
transform 1 0 67804 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_368
timestamp 1649977179
transform 1 0 34960 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_380
timestamp 1649977179
transform 1 0 36064 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1649977179
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1649977179
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1649977179
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1649977179
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1649977179
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1649977179
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1649977179
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1649977179
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1649977179
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1649977179
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1649977179
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_729
timestamp 1649977179
transform 1 0 68172 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1649977179
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1649977179
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1649977179
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1649977179
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1649977179
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1649977179
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1649977179
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1649977179
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1649977179
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1649977179
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1649977179
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1649977179
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1649977179
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_725
timestamp 1649977179
transform 1 0 67804 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1649977179
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1649977179
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1649977179
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1649977179
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1649977179
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1649977179
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1649977179
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1649977179
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1649977179
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1649977179
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1649977179
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1649977179
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_729
timestamp 1649977179
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_64
timestamp 1649977179
transform 1 0 6992 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_76
timestamp 1649977179
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_292
timestamp 1649977179
transform 1 0 27968 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1649977179
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1649977179
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1649977179
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1649977179
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1649977179
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1649977179
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1649977179
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1649977179
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1649977179
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1649977179
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1649977179
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1649977179
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_725
timestamp 1649977179
transform 1 0 67804 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_89
timestamp 1649977179
transform 1 0 9292 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_94
timestamp 1649977179
transform 1 0 9752 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_101
timestamp 1649977179
transform 1 0 10396 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1649977179
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1649977179
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1649977179
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_269
timestamp 1649977179
transform 1 0 25852 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1649977179
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_284
timestamp 1649977179
transform 1 0 27232 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_296
timestamp 1649977179
transform 1 0 28336 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_308
timestamp 1649977179
transform 1 0 29440 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_320
timestamp 1649977179
transform 1 0 30544 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1649977179
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_584
timestamp 1649977179
transform 1 0 54832 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_596
timestamp 1649977179
transform 1 0 55936 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_608
timestamp 1649977179
transform 1 0 57040 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1649977179
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1649977179
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1649977179
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1649977179
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1649977179
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1649977179
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1649977179
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1649977179
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1649977179
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1649977179
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1649977179
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_729
timestamp 1649977179
transform 1 0 68172 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_37
timestamp 1649977179
transform 1 0 4508 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_43
timestamp 1649977179
transform 1 0 5060 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_50
timestamp 1649977179
transform 1 0 5704 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_62
timestamp 1649977179
transform 1 0 6808 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_74
timestamp 1649977179
transform 1 0 7912 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1649977179
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_128
timestamp 1649977179
transform 1 0 12880 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1649977179
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1649977179
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_464
timestamp 1649977179
transform 1 0 43792 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_580
timestamp 1649977179
transform 1 0 54464 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_610
timestamp 1649977179
transform 1 0 57224 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_622
timestamp 1649977179
transform 1 0 58328 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_634
timestamp 1649977179
transform 1 0 59432 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_642
timestamp 1649977179
transform 1 0 60168 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1649977179
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1649977179
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1649977179
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1649977179
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1649977179
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1649977179
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1649977179
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1649977179
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_725
timestamp 1649977179
transform 1 0 67804 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_60
timestamp 1649977179
transform 1 0 6624 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_72
timestamp 1649977179
transform 1 0 7728 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_84
timestamp 1649977179
transform 1 0 8832 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_96
timestamp 1649977179
transform 1 0 9936 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1649977179
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_119
timestamp 1649977179
transform 1 0 12052 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_141
timestamp 1649977179
transform 1 0 14076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_153
timestamp 1649977179
transform 1 0 15180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1649977179
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1649977179
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1649977179
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1649977179
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_483
timestamp 1649977179
transform 1 0 45540 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_495
timestamp 1649977179
transform 1 0 46644 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1649977179
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1649977179
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1649977179
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1649977179
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1649977179
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1649977179
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1649977179
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1649977179
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1649977179
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1649977179
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1649977179
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_729
timestamp 1649977179
transform 1 0 68172 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_45
timestamp 1649977179
transform 1 0 5244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_70
timestamp 1649977179
transform 1 0 7544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_74
timestamp 1649977179
transform 1 0 7912 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_78
timestamp 1649977179
transform 1 0 8280 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_88
timestamp 1649977179
transform 1 0 9200 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_100
timestamp 1649977179
transform 1 0 10304 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_112
timestamp 1649977179
transform 1 0 11408 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_120
timestamp 1649977179
transform 1 0 12144 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_124
timestamp 1649977179
transform 1 0 12512 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1649977179
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1649977179
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1649977179
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1649977179
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1649977179
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1649977179
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_466
timestamp 1649977179
transform 1 0 43976 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_474
timestamp 1649977179
transform 1 0 44712 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1649977179
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1649977179
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1649977179
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1649977179
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1649977179
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1649977179
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1649977179
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1649977179
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1649977179
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1649977179
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_713
timestamp 1649977179
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_725
timestamp 1649977179
transform 1 0 67804 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_96
timestamp 1649977179
transform 1 0 9936 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1649977179
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_285
timestamp 1649977179
transform 1 0 27324 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_297
timestamp 1649977179
transform 1 0 28428 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_309
timestamp 1649977179
transform 1 0 29532 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_321
timestamp 1649977179
transform 1 0 30636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1649977179
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1649977179
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1649977179
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1649977179
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_459
timestamp 1649977179
transform 1 0 43332 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_471
timestamp 1649977179
transform 1 0 44436 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_483
timestamp 1649977179
transform 1 0 45540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_495
timestamp 1649977179
transform 1 0 46644 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1649977179
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1649977179
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1649977179
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1649977179
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1649977179
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1649977179
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1649977179
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1649977179
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1649977179
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1649977179
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1649977179
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_729
timestamp 1649977179
transform 1 0 68172 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_273
timestamp 1649977179
transform 1 0 26220 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_278
timestamp 1649977179
transform 1 0 26680 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1649977179
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1649977179
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_454
timestamp 1649977179
transform 1 0 42872 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_466
timestamp 1649977179
transform 1 0 43976 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_474
timestamp 1649977179
transform 1 0 44712 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_625
timestamp 1649977179
transform 1 0 58604 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_633
timestamp 1649977179
transform 1 0 59340 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_639
timestamp 1649977179
transform 1 0 59892 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1649977179
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1649977179
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1649977179
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1649977179
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1649977179
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1649977179
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1649977179
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1649977179
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1649977179
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_725
timestamp 1649977179
transform 1 0 67804 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_444
timestamp 1649977179
transform 1 0 41952 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_470
timestamp 1649977179
transform 1 0 44344 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_482
timestamp 1649977179
transform 1 0 45448 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_494
timestamp 1649977179
transform 1 0 46552 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_502
timestamp 1649977179
transform 1 0 47288 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_632
timestamp 1649977179
transform 1 0 59248 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_657
timestamp 1649977179
transform 1 0 61548 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_669
timestamp 1649977179
transform 1 0 62652 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1649977179
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1649977179
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1649977179
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1649977179
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_724
timestamp 1649977179
transform 1 0 67712 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_729
timestamp 1649977179
transform 1 0 68172 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1649977179
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_451
timestamp 1649977179
transform 1 0 42596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_463
timestamp 1649977179
transform 1 0 43700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_625
timestamp 1649977179
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1649977179
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1649977179
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1649977179
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1649977179
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1649977179
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1649977179
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1649977179
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1649977179
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_701
timestamp 1649977179
transform 1 0 65596 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_707
timestamp 1649977179
transform 1 0 66148 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_729
timestamp 1649977179
transform 1 0 68172 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1649977179
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_455
timestamp 1649977179
transform 1 0 42964 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_463
timestamp 1649977179
transform 1 0 43700 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_486
timestamp 1649977179
transform 1 0 45816 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_498
timestamp 1649977179
transform 1 0 46920 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1649977179
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1649977179
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_653
timestamp 1649977179
transform 1 0 61180 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_659
timestamp 1649977179
transform 1 0 61732 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_663
timestamp 1649977179
transform 1 0 62100 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1649977179
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1649977179
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1649977179
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_697
timestamp 1649977179
transform 1 0 65228 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_724
timestamp 1649977179
transform 1 0 67712 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_729
timestamp 1649977179
transform 1 0 68172 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1649977179
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_456
timestamp 1649977179
transform 1 0 43056 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_463
timestamp 1649977179
transform 1 0 43700 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_470
timestamp 1649977179
transform 1 0 44344 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1649977179
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1649977179
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1649977179
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1649977179
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_657
timestamp 1649977179
transform 1 0 61548 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_663
timestamp 1649977179
transform 1 0 62100 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_685
timestamp 1649977179
transform 1 0 64124 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_697
timestamp 1649977179
transform 1 0 65228 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1649977179
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_713
timestamp 1649977179
transform 1 0 66700 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_720
timestamp 1649977179
transform 1 0 67344 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_727
timestamp 1649977179
transform 1 0 67988 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_437
timestamp 1649977179
transform 1 0 41308 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_444
timestamp 1649977179
transform 1 0 41952 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_453
timestamp 1649977179
transform 1 0 42780 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_475
timestamp 1649977179
transform 1 0 44804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_487
timestamp 1649977179
transform 1 0 45908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_499
timestamp 1649977179
transform 1 0 47012 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1649977179
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1649977179
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_653
timestamp 1649977179
transform 1 0 61180 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_661
timestamp 1649977179
transform 1 0 61916 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_667
timestamp 1649977179
transform 1 0 62468 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1649977179
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1649977179
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1649977179
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_697
timestamp 1649977179
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_709
timestamp 1649977179
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_724
timestamp 1649977179
transform 1 0 67712 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_729
timestamp 1649977179
transform 1 0 68172 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1649977179
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_455
timestamp 1649977179
transform 1 0 42964 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_462
timestamp 1649977179
transform 1 0 43608 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_474
timestamp 1649977179
transform 1 0 44712 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1649977179
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1649977179
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1649977179
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1649977179
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1649977179
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1649977179
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1649977179
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1649977179
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1649977179
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_701
timestamp 1649977179
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_713
timestamp 1649977179
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_725
timestamp 1649977179
transform 1 0 67804 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1649977179
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1649977179
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1649977179
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1649977179
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1649977179
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1649977179
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_685
timestamp 1649977179
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_697
timestamp 1649977179
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_709
timestamp 1649977179
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1649977179
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1649977179
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_729
timestamp 1649977179
transform 1 0 68172 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_381
timestamp 1649977179
transform 1 0 36156 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_385
timestamp 1649977179
transform 1 0 36524 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_410
timestamp 1649977179
transform 1 0 38824 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_418
timestamp 1649977179
transform 1 0 39560 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_625
timestamp 1649977179
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1649977179
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1649977179
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_645
timestamp 1649977179
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_657
timestamp 1649977179
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_669
timestamp 1649977179
transform 1 0 62652 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_676
timestamp 1649977179
transform 1 0 63296 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_683
timestamp 1649977179
transform 1 0 63940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_695
timestamp 1649977179
transform 1 0 65044 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1649977179
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_701
timestamp 1649977179
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_713
timestamp 1649977179
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_725
timestamp 1649977179
transform 1 0 67804 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_397
timestamp 1649977179
transform 1 0 37628 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_401
timestamp 1649977179
transform 1 0 37996 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_423
timestamp 1649977179
transform 1 0 40020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_435
timestamp 1649977179
transform 1 0 41124 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_629
timestamp 1649977179
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_641
timestamp 1649977179
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_653
timestamp 1649977179
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1649977179
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1649977179
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_694
timestamp 1649977179
transform 1 0 64952 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_706
timestamp 1649977179
transform 1 0 66056 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_718
timestamp 1649977179
transform 1 0 67160 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_726
timestamp 1649977179
transform 1 0 67896 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_729
timestamp 1649977179
transform 1 0 68172 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_66
timestamp 1649977179
transform 1 0 7176 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_78
timestamp 1649977179
transform 1 0 8280 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_214
timestamp 1649977179
transform 1 0 20792 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_226
timestamp 1649977179
transform 1 0 21896 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_238
timestamp 1649977179
transform 1 0 23000 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1649977179
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1649977179
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1649977179
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1649977179
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_625
timestamp 1649977179
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1649977179
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1649977179
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_645
timestamp 1649977179
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_657
timestamp 1649977179
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_669
timestamp 1649977179
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_681
timestamp 1649977179
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1649977179
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1649977179
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_701
timestamp 1649977179
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_713
timestamp 1649977179
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_725
timestamp 1649977179
transform 1 0 67804 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_50
timestamp 1649977179
transform 1 0 5704 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_78
timestamp 1649977179
transform 1 0 8280 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_90
timestamp 1649977179
transform 1 0 9384 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_102
timestamp 1649977179
transform 1 0 10488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1649977179
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_211
timestamp 1649977179
transform 1 0 20516 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_218
timestamp 1649977179
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_401
timestamp 1649977179
transform 1 0 37996 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_406
timestamp 1649977179
transform 1 0 38456 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_413
timestamp 1649977179
transform 1 0 39100 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_425
timestamp 1649977179
transform 1 0 40204 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_437
timestamp 1649977179
transform 1 0 41308 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_445
timestamp 1649977179
transform 1 0 42044 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_629
timestamp 1649977179
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_641
timestamp 1649977179
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_653
timestamp 1649977179
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1649977179
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1649977179
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_673
timestamp 1649977179
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_685
timestamp 1649977179
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_697
timestamp 1649977179
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_709
timestamp 1649977179
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1649977179
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1649977179
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_729
timestamp 1649977179
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1649977179
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_59
timestamp 1649977179
transform 1 0 6532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_71
timestamp 1649977179
transform 1 0 7636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_201
timestamp 1649977179
transform 1 0 19596 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_208
timestamp 1649977179
transform 1 0 20240 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_218
timestamp 1649977179
transform 1 0 21160 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_228
timestamp 1649977179
transform 1 0 22080 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_240
timestamp 1649977179
transform 1 0 23184 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1649977179
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1649977179
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1649977179
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_567
timestamp 1649977179
transform 1 0 53268 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_579
timestamp 1649977179
transform 1 0 54372 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_625
timestamp 1649977179
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_637
timestamp 1649977179
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1649977179
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_645
timestamp 1649977179
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_657
timestamp 1649977179
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_669
timestamp 1649977179
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_681
timestamp 1649977179
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_693
timestamp 1649977179
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_699
timestamp 1649977179
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_701
timestamp 1649977179
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_713
timestamp 1649977179
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_725
timestamp 1649977179
transform 1 0 67804 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_63
timestamp 1649977179
transform 1 0 6900 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_75
timestamp 1649977179
transform 1 0 8004 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_87
timestamp 1649977179
transform 1 0 9108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_99
timestamp 1649977179
transform 1 0 10212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_236
timestamp 1649977179
transform 1 0 22816 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_248
timestamp 1649977179
transform 1 0 23920 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_260
timestamp 1649977179
transform 1 0 25024 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_272
timestamp 1649977179
transform 1 0 26128 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1649977179
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_343
timestamp 1649977179
transform 1 0 32660 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_347
timestamp 1649977179
transform 1 0 33028 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_354
timestamp 1649977179
transform 1 0 33672 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_366
timestamp 1649977179
transform 1 0 34776 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_378
timestamp 1649977179
transform 1 0 35880 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_390
timestamp 1649977179
transform 1 0 36984 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_524
timestamp 1649977179
transform 1 0 49312 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_536
timestamp 1649977179
transform 1 0 50416 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_547
timestamp 1649977179
transform 1 0 51428 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_629
timestamp 1649977179
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_641
timestamp 1649977179
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_653
timestamp 1649977179
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1649977179
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_671
timestamp 1649977179
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_673
timestamp 1649977179
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_685
timestamp 1649977179
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_697
timestamp 1649977179
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_709
timestamp 1649977179
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_721
timestamp 1649977179
transform 1 0 67436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_727
timestamp 1649977179
transform 1 0 67988 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_729
timestamp 1649977179
transform 1 0 68172 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_217
timestamp 1649977179
transform 1 0 21068 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_223
timestamp 1649977179
transform 1 0 21620 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_248
timestamp 1649977179
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_360
timestamp 1649977179
transform 1 0 34224 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_472
timestamp 1649977179
transform 1 0 44528 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_498
timestamp 1649977179
transform 1 0 46920 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_510
timestamp 1649977179
transform 1 0 48024 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_522
timestamp 1649977179
transform 1 0 49128 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_530
timestamp 1649977179
transform 1 0 49864 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_549
timestamp 1649977179
transform 1 0 51612 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_561
timestamp 1649977179
transform 1 0 52716 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_573
timestamp 1649977179
transform 1 0 53820 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_585
timestamp 1649977179
transform 1 0 54924 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_625
timestamp 1649977179
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_637
timestamp 1649977179
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_643
timestamp 1649977179
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_645
timestamp 1649977179
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_657
timestamp 1649977179
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_669
timestamp 1649977179
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_681
timestamp 1649977179
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_693
timestamp 1649977179
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_699
timestamp 1649977179
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_701
timestamp 1649977179
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_713
timestamp 1649977179
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_725
timestamp 1649977179
transform 1 0 67804 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_97
timestamp 1649977179
transform 1 0 10028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_109
timestamp 1649977179
transform 1 0 11132 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_229
timestamp 1649977179
transform 1 0 22172 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_251
timestamp 1649977179
transform 1 0 24196 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_263
timestamp 1649977179
transform 1 0 25300 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_275
timestamp 1649977179
transform 1 0 26404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1649977179
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_365
timestamp 1649977179
transform 1 0 34684 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_369
timestamp 1649977179
transform 1 0 35052 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_381
timestamp 1649977179
transform 1 0 36156 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_389
timestamp 1649977179
transform 1 0 36892 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_476
timestamp 1649977179
transform 1 0 44896 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_488
timestamp 1649977179
transform 1 0 46000 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_500
timestamp 1649977179
transform 1 0 47104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_512
timestamp 1649977179
transform 1 0 48208 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_524
timestamp 1649977179
transform 1 0 49312 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_536
timestamp 1649977179
transform 1 0 50416 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_548
timestamp 1649977179
transform 1 0 51520 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_629
timestamp 1649977179
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_641
timestamp 1649977179
transform 1 0 60076 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_647
timestamp 1649977179
transform 1 0 60628 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_659
timestamp 1649977179
transform 1 0 61732 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1649977179
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_673
timestamp 1649977179
transform 1 0 63020 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_680
timestamp 1649977179
transform 1 0 63664 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_692
timestamp 1649977179
transform 1 0 64768 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_704
timestamp 1649977179
transform 1 0 65872 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_716
timestamp 1649977179
transform 1 0 66976 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_729
timestamp 1649977179
transform 1 0 68172 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_91
timestamp 1649977179
transform 1 0 9476 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_113
timestamp 1649977179
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_125
timestamp 1649977179
transform 1 0 12604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_137
timestamp 1649977179
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_229
timestamp 1649977179
transform 1 0 22172 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_233
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_240
timestamp 1649977179
transform 1 0 23184 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1649977179
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1649977179
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1649977179
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_390
timestamp 1649977179
transform 1 0 36984 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_402
timestamp 1649977179
transform 1 0 38088 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_414
timestamp 1649977179
transform 1 0 39192 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_625
timestamp 1649977179
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_637
timestamp 1649977179
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1649977179
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_666
timestamp 1649977179
transform 1 0 62376 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_674
timestamp 1649977179
transform 1 0 63112 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_696
timestamp 1649977179
transform 1 0 65136 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_701
timestamp 1649977179
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_713
timestamp 1649977179
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_725
timestamp 1649977179
transform 1 0 67804 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1649977179
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1649977179
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_89
timestamp 1649977179
transform 1 0 9292 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_95
timestamp 1649977179
transform 1 0 9844 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_107
timestamp 1649977179
transform 1 0 10948 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1649977179
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1649977179
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_369
timestamp 1649977179
transform 1 0 35052 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_629
timestamp 1649977179
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_641
timestamp 1649977179
transform 1 0 60076 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_645
timestamp 1649977179
transform 1 0 60444 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_649
timestamp 1649977179
transform 1 0 60812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_661
timestamp 1649977179
transform 1 0 61916 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_669
timestamp 1649977179
transform 1 0 62652 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_673
timestamp 1649977179
transform 1 0 63020 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_679
timestamp 1649977179
transform 1 0 63572 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_683
timestamp 1649977179
transform 1 0 63940 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_695
timestamp 1649977179
transform 1 0 65044 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_707
timestamp 1649977179
transform 1 0 66148 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_719
timestamp 1649977179
transform 1 0 67252 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_727
timestamp 1649977179
transform 1 0 67988 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_729
timestamp 1649977179
transform 1 0 68172 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_618
timestamp 1649977179
transform 1 0 57960 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_630
timestamp 1649977179
transform 1 0 59064 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_642
timestamp 1649977179
transform 1 0 60168 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_645
timestamp 1649977179
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_657
timestamp 1649977179
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_669
timestamp 1649977179
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_681
timestamp 1649977179
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1649977179
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1649977179
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_701
timestamp 1649977179
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_713
timestamp 1649977179
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_725
timestamp 1649977179
transform 1 0 67804 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1649977179
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1649977179
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1649977179
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_612
timestamp 1649977179
transform 1 0 57408 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_638
timestamp 1649977179
transform 1 0 59800 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_650
timestamp 1649977179
transform 1 0 60904 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_662
timestamp 1649977179
transform 1 0 62008 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_670
timestamp 1649977179
transform 1 0 62744 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_673
timestamp 1649977179
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_685
timestamp 1649977179
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_697
timestamp 1649977179
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_709
timestamp 1649977179
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_721
timestamp 1649977179
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_727
timestamp 1649977179
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_729
timestamp 1649977179
transform 1 0 68172 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1649977179
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_625
timestamp 1649977179
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_637
timestamp 1649977179
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1649977179
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_645
timestamp 1649977179
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_657
timestamp 1649977179
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_669
timestamp 1649977179
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_681
timestamp 1649977179
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1649977179
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1649977179
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_701
timestamp 1649977179
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_713
timestamp 1649977179
transform 1 0 66700 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_725
timestamp 1649977179
transform 1 0 67804 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_216
timestamp 1649977179
transform 1 0 20976 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_579
timestamp 1649977179
transform 1 0 54372 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_604
timestamp 1649977179
transform 1 0 56672 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_629
timestamp 1649977179
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_641
timestamp 1649977179
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_653
timestamp 1649977179
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1649977179
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1649977179
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_673
timestamp 1649977179
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_685
timestamp 1649977179
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_697
timestamp 1649977179
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_709
timestamp 1649977179
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_721
timestamp 1649977179
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_727
timestamp 1649977179
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_729
timestamp 1649977179
transform 1 0 68172 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_577
timestamp 1649977179
transform 1 0 54188 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_583
timestamp 1649977179
transform 1 0 54740 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_625
timestamp 1649977179
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_637
timestamp 1649977179
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_643
timestamp 1649977179
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_645
timestamp 1649977179
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_657
timestamp 1649977179
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_669
timestamp 1649977179
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_681
timestamp 1649977179
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1649977179
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1649977179
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_701
timestamp 1649977179
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_713
timestamp 1649977179
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_725
timestamp 1649977179
transform 1 0 67804 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_565
timestamp 1649977179
transform 1 0 53084 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_577
timestamp 1649977179
transform 1 0 54188 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_589
timestamp 1649977179
transform 1 0 55292 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_601
timestamp 1649977179
transform 1 0 56396 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_613
timestamp 1649977179
transform 1 0 57500 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_629
timestamp 1649977179
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_641
timestamp 1649977179
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_653
timestamp 1649977179
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1649977179
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1649977179
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_673
timestamp 1649977179
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_685
timestamp 1649977179
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_697
timestamp 1649977179
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_709
timestamp 1649977179
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_721
timestamp 1649977179
transform 1 0 67436 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_727
timestamp 1649977179
transform 1 0 67988 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_729
timestamp 1649977179
transform 1 0 68172 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_553
timestamp 1649977179
transform 1 0 51980 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_582
timestamp 1649977179
transform 1 0 54648 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_625
timestamp 1649977179
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1649977179
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1649977179
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_645
timestamp 1649977179
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_657
timestamp 1649977179
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_669
timestamp 1649977179
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_681
timestamp 1649977179
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1649977179
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1649977179
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_701
timestamp 1649977179
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_713
timestamp 1649977179
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_725
timestamp 1649977179
transform 1 0 67804 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_154
timestamp 1649977179
transform 1 0 15272 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_166
timestamp 1649977179
transform 1 0 16376 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_397
timestamp 1649977179
transform 1 0 37628 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_404
timestamp 1649977179
transform 1 0 38272 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_416
timestamp 1649977179
transform 1 0 39376 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_428
timestamp 1649977179
transform 1 0 40480 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_440
timestamp 1649977179
transform 1 0 41584 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_465
timestamp 1649977179
transform 1 0 43884 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_470
timestamp 1649977179
transform 1 0 44344 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_482
timestamp 1649977179
transform 1 0 45448 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_494
timestamp 1649977179
transform 1 0 46552 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_502
timestamp 1649977179
transform 1 0 47288 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_629
timestamp 1649977179
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_641
timestamp 1649977179
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_653
timestamp 1649977179
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1649977179
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1649977179
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_673
timestamp 1649977179
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_685
timestamp 1649977179
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_697
timestamp 1649977179
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_709
timestamp 1649977179
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_724
timestamp 1649977179
transform 1 0 67712 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_729
timestamp 1649977179
transform 1 0 68172 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_147
timestamp 1649977179
transform 1 0 14628 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_169
timestamp 1649977179
transform 1 0 16652 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_181
timestamp 1649977179
transform 1 0 17756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_193
timestamp 1649977179
transform 1 0 18860 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_385
timestamp 1649977179
transform 1 0 36524 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_391
timestamp 1649977179
transform 1 0 37076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_403
timestamp 1649977179
transform 1 0 38180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_415
timestamp 1649977179
transform 1 0 39284 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_625
timestamp 1649977179
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1649977179
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1649977179
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_645
timestamp 1649977179
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_657
timestamp 1649977179
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_669
timestamp 1649977179
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_681
timestamp 1649977179
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1649977179
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1649977179
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_701
timestamp 1649977179
transform 1 0 65596 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_707
timestamp 1649977179
transform 1 0 66148 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_729
timestamp 1649977179
transform 1 0 68172 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_145
timestamp 1649977179
transform 1 0 14444 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_151
timestamp 1649977179
transform 1 0 14996 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_163
timestamp 1649977179
transform 1 0 16100 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_414
timestamp 1649977179
transform 1 0 39192 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_426
timestamp 1649977179
transform 1 0 40296 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_438
timestamp 1649977179
transform 1 0 41400 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_446
timestamp 1649977179
transform 1 0 42136 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_531
timestamp 1649977179
transform 1 0 49956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_543
timestamp 1649977179
transform 1 0 51060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_555
timestamp 1649977179
transform 1 0 52164 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_629
timestamp 1649977179
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_641
timestamp 1649977179
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_653
timestamp 1649977179
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1649977179
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1649977179
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_673
timestamp 1649977179
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_685
timestamp 1649977179
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_697
timestamp 1649977179
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_709
timestamp 1649977179
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_724
timestamp 1649977179
transform 1 0 67712 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_729
timestamp 1649977179
transform 1 0 68172 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_395
timestamp 1649977179
transform 1 0 37444 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_407
timestamp 1649977179
transform 1 0 38548 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_625
timestamp 1649977179
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1649977179
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1649977179
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_645
timestamp 1649977179
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_657
timestamp 1649977179
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_669
timestamp 1649977179
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_681
timestamp 1649977179
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_693
timestamp 1649977179
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_699
timestamp 1649977179
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_701
timestamp 1649977179
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_713
timestamp 1649977179
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_725
timestamp 1649977179
transform 1 0 67804 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_629
timestamp 1649977179
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_641
timestamp 1649977179
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_653
timestamp 1649977179
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_665
timestamp 1649977179
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_671
timestamp 1649977179
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_673
timestamp 1649977179
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_685
timestamp 1649977179
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_697
timestamp 1649977179
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_709
timestamp 1649977179
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_721
timestamp 1649977179
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_727
timestamp 1649977179
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_729
timestamp 1649977179
transform 1 0 68172 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_461
timestamp 1649977179
transform 1 0 43516 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1649977179
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_486
timestamp 1649977179
transform 1 0 45816 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_498
timestamp 1649977179
transform 1 0 46920 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_510
timestamp 1649977179
transform 1 0 48024 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_522
timestamp 1649977179
transform 1 0 49128 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_530
timestamp 1649977179
transform 1 0 49864 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_625
timestamp 1649977179
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_637
timestamp 1649977179
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_643
timestamp 1649977179
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_645
timestamp 1649977179
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_657
timestamp 1649977179
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_669
timestamp 1649977179
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_681
timestamp 1649977179
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_693
timestamp 1649977179
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_699
timestamp 1649977179
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_704
timestamp 1649977179
transform 1 0 65872 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_716
timestamp 1649977179
transform 1 0 66976 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_728
timestamp 1649977179
transform 1 0 68080 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_732
timestamp 1649977179
transform 1 0 68448 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_457
timestamp 1649977179
transform 1 0 43148 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_481
timestamp 1649977179
transform 1 0 45356 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_493
timestamp 1649977179
transform 1 0 46460 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_501
timestamp 1649977179
transform 1 0 47196 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_629
timestamp 1649977179
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_641
timestamp 1649977179
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_653
timestamp 1649977179
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_665
timestamp 1649977179
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_671
timestamp 1649977179
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_673
timestamp 1649977179
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_685
timestamp 1649977179
transform 1 0 64124 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_694
timestamp 1649977179
transform 1 0 64952 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_719
timestamp 1649977179
transform 1 0 67252 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_727
timestamp 1649977179
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_729
timestamp 1649977179
transform 1 0 68172 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1649977179
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1649977179
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1649977179
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_453
timestamp 1649977179
transform 1 0 42780 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_459
timestamp 1649977179
transform 1 0 43332 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_483
timestamp 1649977179
transform 1 0 45540 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_495
timestamp 1649977179
transform 1 0 46644 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_507
timestamp 1649977179
transform 1 0 47748 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_519
timestamp 1649977179
transform 1 0 48852 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_625
timestamp 1649977179
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1649977179
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1649977179
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_645
timestamp 1649977179
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_657
timestamp 1649977179
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_669
timestamp 1649977179
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_681
timestamp 1649977179
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1649977179
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1649977179
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_701
timestamp 1649977179
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_713
timestamp 1649977179
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_725
timestamp 1649977179
transform 1 0 67804 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_464
timestamp 1649977179
transform 1 0 43792 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_474
timestamp 1649977179
transform 1 0 44712 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_484
timestamp 1649977179
transform 1 0 45632 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_496
timestamp 1649977179
transform 1 0 46736 0 -1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_565
timestamp 1649977179
transform 1 0 53084 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_569
timestamp 1649977179
transform 1 0 53452 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_594
timestamp 1649977179
transform 1 0 55752 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_606
timestamp 1649977179
transform 1 0 56856 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_614
timestamp 1649977179
transform 1 0 57592 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_629
timestamp 1649977179
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_641
timestamp 1649977179
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_653
timestamp 1649977179
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1649977179
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1649977179
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_673
timestamp 1649977179
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_685
timestamp 1649977179
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_697
timestamp 1649977179
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_709
timestamp 1649977179
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_721
timestamp 1649977179
transform 1 0 67436 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_727
timestamp 1649977179
transform 1 0 67988 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_729
timestamp 1649977179
transform 1 0 68172 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1649977179
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_69
timestamp 1649977179
transform 1 0 7452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_81
timestamp 1649977179
transform 1 0 8556 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_297
timestamp 1649977179
transform 1 0 28428 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_86_320
timestamp 1649977179
transform 1 0 30544 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_332
timestamp 1649977179
transform 1 0 31648 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_344
timestamp 1649977179
transform 1 0 32752 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_356
timestamp 1649977179
transform 1 0 33856 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_573
timestamp 1649977179
transform 1 0 53820 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_577
timestamp 1649977179
transform 1 0 54188 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_585
timestamp 1649977179
transform 1 0 54924 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_625
timestamp 1649977179
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1649977179
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1649977179
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_645
timestamp 1649977179
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_657
timestamp 1649977179
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_669
timestamp 1649977179
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_681
timestamp 1649977179
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1649977179
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1649977179
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_701
timestamp 1649977179
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_713
timestamp 1649977179
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_725
timestamp 1649977179
transform 1 0 67804 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_84
timestamp 1649977179
transform 1 0 8832 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_96
timestamp 1649977179
transform 1 0 9936 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_108
timestamp 1649977179
transform 1 0 11040 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_285
timestamp 1649977179
transform 1 0 27324 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_307
timestamp 1649977179
transform 1 0 29348 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_332
timestamp 1649977179
transform 1 0 31648 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1649977179
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1649977179
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1649977179
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_629
timestamp 1649977179
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_641
timestamp 1649977179
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_653
timestamp 1649977179
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1649977179
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1649977179
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_673
timestamp 1649977179
transform 1 0 63020 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_677
timestamp 1649977179
transform 1 0 63388 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_689
timestamp 1649977179
transform 1 0 64492 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_701
timestamp 1649977179
transform 1 0 65596 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_713
timestamp 1649977179
transform 1 0 66700 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_725
timestamp 1649977179
transform 1 0 67804 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_729
timestamp 1649977179
transform 1 0 68172 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1649977179
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1649977179
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1649977179
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_61
timestamp 1649977179
transform 1 0 6716 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_67
timestamp 1649977179
transform 1 0 7268 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_79
timestamp 1649977179
transform 1 0 8372 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_297
timestamp 1649977179
transform 1 0 28428 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_318
timestamp 1649977179
transform 1 0 30360 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_330
timestamp 1649977179
transform 1 0 31464 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_342
timestamp 1649977179
transform 1 0 32568 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_354
timestamp 1649977179
transform 1 0 33672 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_362
timestamp 1649977179
transform 1 0 34408 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_374
timestamp 1649977179
transform 1 0 35512 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_386
timestamp 1649977179
transform 1 0 36616 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_398
timestamp 1649977179
transform 1 0 37720 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_410
timestamp 1649977179
transform 1 0 38824 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_418
timestamp 1649977179
transform 1 0 39560 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_485
timestamp 1649977179
transform 1 0 45724 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_490
timestamp 1649977179
transform 1 0 46184 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_502
timestamp 1649977179
transform 1 0 47288 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_514
timestamp 1649977179
transform 1 0 48392 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_526
timestamp 1649977179
transform 1 0 49496 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1649977179
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1649977179
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_625
timestamp 1649977179
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1649977179
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1649977179
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_645
timestamp 1649977179
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_657
timestamp 1649977179
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_669
timestamp 1649977179
transform 1 0 62652 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_88_696
timestamp 1649977179
transform 1 0 65136 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_701
timestamp 1649977179
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_713
timestamp 1649977179
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_725
timestamp 1649977179
transform 1 0 67804 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1649977179
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1649977179
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1649977179
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1649977179
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_89_388
timestamp 1649977179
transform 1 0 36800 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_89_500
timestamp 1649977179
transform 1 0 47104 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_548
timestamp 1649977179
transform 1 0 51520 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1649977179
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1649977179
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1649977179
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1649977179
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1649977179
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_629
timestamp 1649977179
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_641
timestamp 1649977179
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_653
timestamp 1649977179
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1649977179
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1649977179
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_673
timestamp 1649977179
transform 1 0 63020 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_677
timestamp 1649977179
transform 1 0 63388 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_681
timestamp 1649977179
transform 1 0 63756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_693
timestamp 1649977179
transform 1 0 64860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_705
timestamp 1649977179
transform 1 0 65964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_717
timestamp 1649977179
transform 1 0 67068 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_725
timestamp 1649977179
transform 1 0 67804 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_729
timestamp 1649977179
transform 1 0 68172 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1649977179
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1649977179
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_371
timestamp 1649977179
transform 1 0 35236 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_375
timestamp 1649977179
transform 1 0 35604 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_387
timestamp 1649977179
transform 1 0 36708 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_399
timestamp 1649977179
transform 1 0 37812 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_411
timestamp 1649977179
transform 1 0 38916 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_484
timestamp 1649977179
transform 1 0 45632 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_496
timestamp 1649977179
transform 1 0 46736 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_508
timestamp 1649977179
transform 1 0 47840 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_520
timestamp 1649977179
transform 1 0 48944 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_567
timestamp 1649977179
transform 1 0 53268 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_579
timestamp 1649977179
transform 1 0 54372 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_625
timestamp 1649977179
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1649977179
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1649977179
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_645
timestamp 1649977179
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_657
timestamp 1649977179
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_669
timestamp 1649977179
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_681
timestamp 1649977179
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1649977179
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1649977179
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_701
timestamp 1649977179
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_713
timestamp 1649977179
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_725
timestamp 1649977179
transform 1 0 67804 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1649977179
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1649977179
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_39
timestamp 1649977179
transform 1 0 4692 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_47
timestamp 1649977179
transform 1 0 5428 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_52
timestamp 1649977179
transform 1 0 5888 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_91
timestamp 1649977179
transform 1 0 9476 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_103
timestamp 1649977179
transform 1 0 10580 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_91_550
timestamp 1649977179
transform 1 0 51704 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_558
timestamp 1649977179
transform 1 0 52440 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1649977179
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1649977179
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1649977179
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1649977179
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_629
timestamp 1649977179
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_641
timestamp 1649977179
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_653
timestamp 1649977179
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1649977179
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1649977179
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_673
timestamp 1649977179
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_685
timestamp 1649977179
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_697
timestamp 1649977179
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_709
timestamp 1649977179
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_721
timestamp 1649977179
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_727
timestamp 1649977179
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_729
timestamp 1649977179
transform 1 0 68172 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1649977179
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1649977179
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1649977179
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_66
timestamp 1649977179
transform 1 0 7176 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_74
timestamp 1649977179
transform 1 0 7912 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_79
timestamp 1649977179
transform 1 0 8372 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1649977179
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1649977179
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_625
timestamp 1649977179
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1649977179
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1649977179
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_645
timestamp 1649977179
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_657
timestamp 1649977179
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_669
timestamp 1649977179
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_681
timestamp 1649977179
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1649977179
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1649977179
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_701
timestamp 1649977179
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_713
timestamp 1649977179
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_725
timestamp 1649977179
transform 1 0 67804 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1649977179
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1649977179
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_39
timestamp 1649977179
transform 1 0 4692 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_45
timestamp 1649977179
transform 1 0 5244 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_49
timestamp 1649977179
transform 1 0 5612 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_74
timestamp 1649977179
transform 1 0 7912 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_86
timestamp 1649977179
transform 1 0 9016 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_98
timestamp 1649977179
transform 1 0 10120 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1649977179
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_289
timestamp 1649977179
transform 1 0 27692 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_401
timestamp 1649977179
transform 1 0 37996 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_406
timestamp 1649977179
transform 1 0 38456 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_431
timestamp 1649977179
transform 1 0 40756 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_443
timestamp 1649977179
transform 1 0 41860 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_546
timestamp 1649977179
transform 1 0 51336 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_558
timestamp 1649977179
transform 1 0 52440 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1649977179
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1649977179
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1649977179
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1649977179
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1649977179
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_629
timestamp 1649977179
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_641
timestamp 1649977179
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_653
timestamp 1649977179
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1649977179
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1649977179
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_673
timestamp 1649977179
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_685
timestamp 1649977179
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_697
timestamp 1649977179
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_709
timestamp 1649977179
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_724
timestamp 1649977179
transform 1 0 67712 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_729
timestamp 1649977179
transform 1 0 68172 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1649977179
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1649977179
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_94_304
timestamp 1649977179
transform 1 0 29072 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_541
timestamp 1649977179
transform 1 0 50876 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_565
timestamp 1649977179
transform 1 0 53084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_577
timestamp 1649977179
transform 1 0 54188 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_585
timestamp 1649977179
transform 1 0 54924 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_625
timestamp 1649977179
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1649977179
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1649977179
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_645
timestamp 1649977179
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_657
timestamp 1649977179
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_669
timestamp 1649977179
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_681
timestamp 1649977179
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1649977179
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1649977179
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_701
timestamp 1649977179
transform 1 0 65596 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_707
timestamp 1649977179
transform 1 0 66148 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_729
timestamp 1649977179
transform 1 0 68172 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1649977179
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1649977179
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1649977179
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1649977179
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_288
timestamp 1649977179
transform 1 0 27600 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_300
timestamp 1649977179
transform 1 0 28704 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_312
timestamp 1649977179
transform 1 0 29808 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_324
timestamp 1649977179
transform 1 0 30912 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_409
timestamp 1649977179
transform 1 0 38732 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_413
timestamp 1649977179
transform 1 0 39100 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_425
timestamp 1649977179
transform 1 0 40204 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_437
timestamp 1649977179
transform 1 0 41308 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_445
timestamp 1649977179
transform 1 0 42044 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_548
timestamp 1649977179
transform 1 0 51520 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1649977179
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_629
timestamp 1649977179
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_641
timestamp 1649977179
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_653
timestamp 1649977179
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1649977179
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1649977179
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_673
timestamp 1649977179
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_685
timestamp 1649977179
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_697
timestamp 1649977179
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_709
timestamp 1649977179
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_724
timestamp 1649977179
transform 1 0 67712 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_729
timestamp 1649977179
transform 1 0 68172 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1649977179
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1649977179
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1649977179
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_625
timestamp 1649977179
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_637
timestamp 1649977179
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_643
timestamp 1649977179
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_645
timestamp 1649977179
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_657
timestamp 1649977179
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_669
timestamp 1649977179
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_681
timestamp 1649977179
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_693
timestamp 1649977179
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_699
timestamp 1649977179
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_701
timestamp 1649977179
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_713
timestamp 1649977179
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_725
timestamp 1649977179
transform 1 0 67804 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1649977179
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1649977179
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1649977179
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1649977179
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1649977179
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1649977179
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1649977179
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1649977179
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1649977179
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1649977179
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1649977179
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_341
timestamp 1649977179
transform 1 0 32476 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_363
timestamp 1649977179
transform 1 0 34500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_375
timestamp 1649977179
transform 1 0 35604 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_387
timestamp 1649977179
transform 1 0 36708 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_396
timestamp 1649977179
transform 1 0 37536 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_408
timestamp 1649977179
transform 1 0 38640 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_420
timestamp 1649977179
transform 1 0 39744 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_432
timestamp 1649977179
transform 1 0 40848 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_444
timestamp 1649977179
transform 1 0 41952 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_597
timestamp 1649977179
transform 1 0 56028 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_605
timestamp 1649977179
transform 1 0 56764 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_97_610
timestamp 1649977179
transform 1 0 57224 0 -1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_638
timestamp 1649977179
transform 1 0 59800 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_650
timestamp 1649977179
transform 1 0 60904 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_662
timestamp 1649977179
transform 1 0 62008 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_670
timestamp 1649977179
transform 1 0 62744 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_673
timestamp 1649977179
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_685
timestamp 1649977179
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_697
timestamp 1649977179
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_709
timestamp 1649977179
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_721
timestamp 1649977179
transform 1 0 67436 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_727
timestamp 1649977179
transform 1 0 67988 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_729
timestamp 1649977179
transform 1 0 68172 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1649977179
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1649977179
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1649977179
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1649977179
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1649977179
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1649977179
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1649977179
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1649977179
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1649977179
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1649977179
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1649977179
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1649977179
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1649977179
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1649977179
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1649977179
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1649977179
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1649977179
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1649977179
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1649977179
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1649977179
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1649977179
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1649977179
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1649977179
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1649977179
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1649977179
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1649977179
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1649977179
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1649977179
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1649977179
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1649977179
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1649977179
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1649977179
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_601
timestamp 1649977179
transform 1 0 56396 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_98_612
timestamp 1649977179
transform 1 0 57408 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_624
timestamp 1649977179
transform 1 0 58512 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_636
timestamp 1649977179
transform 1 0 59616 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_98_645
timestamp 1649977179
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_657
timestamp 1649977179
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_669
timestamp 1649977179
transform 1 0 62652 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_681
timestamp 1649977179
transform 1 0 63756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_693
timestamp 1649977179
transform 1 0 64860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_699
timestamp 1649977179
transform 1 0 65412 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_701
timestamp 1649977179
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_713
timestamp 1649977179
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_725
timestamp 1649977179
transform 1 0 67804 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1649977179
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1649977179
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1649977179
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1649977179
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_116
timestamp 1649977179
transform 1 0 11776 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_128
timestamp 1649977179
transform 1 0 12880 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_140
timestamp 1649977179
transform 1 0 13984 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_152
timestamp 1649977179
transform 1 0 15088 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_164
timestamp 1649977179
transform 1 0 16192 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1649977179
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1649977179
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1649977179
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1649977179
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1649977179
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1649977179
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1649977179
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1649977179
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1649977179
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1649977179
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1649977179
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1649977179
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1649977179
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1649977179
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1649977179
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1649977179
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1649977179
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1649977179
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1649977179
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1649977179
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1649977179
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1649977179
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1649977179
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1649977179
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1649977179
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1649977179
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1649977179
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1649977179
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_617
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_629
timestamp 1649977179
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_641
timestamp 1649977179
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_653
timestamp 1649977179
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_665
timestamp 1649977179
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1649977179
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_673
timestamp 1649977179
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_685
timestamp 1649977179
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_697
timestamp 1649977179
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_709
timestamp 1649977179
transform 1 0 66332 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_721
timestamp 1649977179
transform 1 0 67436 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_727
timestamp 1649977179
transform 1 0 67988 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_729
timestamp 1649977179
transform 1 0 68172 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1649977179
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1649977179
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1649977179
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_101
timestamp 1649977179
transform 1 0 10396 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_105
timestamp 1649977179
transform 1 0 10764 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_130
timestamp 1649977179
transform 1 0 13064 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_138
timestamp 1649977179
transform 1 0 13800 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1649977179
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1649977179
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1649977179
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1649977179
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1649977179
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1649977179
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1649977179
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1649977179
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1649977179
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1649977179
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1649977179
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1649977179
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1649977179
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1649977179
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1649977179
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1649977179
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1649977179
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1649977179
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1649977179
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1649977179
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1649977179
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1649977179
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1649977179
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1649977179
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1649977179
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1649977179
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1649977179
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1649977179
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_513
timestamp 1649977179
transform 1 0 48300 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_518
timestamp 1649977179
transform 1 0 48760 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_530
timestamp 1649977179
transform 1 0 49864 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1649977179
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_625
timestamp 1649977179
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_637
timestamp 1649977179
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_643
timestamp 1649977179
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_645
timestamp 1649977179
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_657
timestamp 1649977179
transform 1 0 61548 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_669
timestamp 1649977179
transform 1 0 62652 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_681
timestamp 1649977179
transform 1 0 63756 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_693
timestamp 1649977179
transform 1 0 64860 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_699
timestamp 1649977179
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_701
timestamp 1649977179
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_713
timestamp 1649977179
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_725
timestamp 1649977179
transform 1 0 67804 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1649977179
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_27
timestamp 1649977179
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_39
timestamp 1649977179
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1649977179
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1649977179
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1649977179
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_81
timestamp 1649977179
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_93
timestamp 1649977179
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1649977179
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1649977179
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1649977179
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1649977179
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_137
timestamp 1649977179
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_149
timestamp 1649977179
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_161
timestamp 1649977179
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1649977179
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1649977179
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1649977179
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_193
timestamp 1649977179
transform 1 0 18860 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_205
timestamp 1649977179
transform 1 0 19964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_217
timestamp 1649977179
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1649977179
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1649977179
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1649977179
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_249
timestamp 1649977179
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_261
timestamp 1649977179
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1649977179
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1649977179
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1649977179
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1649977179
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_305
timestamp 1649977179
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_317
timestamp 1649977179
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_329
timestamp 1649977179
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_335
timestamp 1649977179
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1649977179
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1649977179
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_361
timestamp 1649977179
transform 1 0 34316 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_373
timestamp 1649977179
transform 1 0 35420 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_385
timestamp 1649977179
transform 1 0 36524 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_391
timestamp 1649977179
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1649977179
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1649977179
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_417
timestamp 1649977179
transform 1 0 39468 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_429
timestamp 1649977179
transform 1 0 40572 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1649977179
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1649977179
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1649977179
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1649977179
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_473
timestamp 1649977179
transform 1 0 44620 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_485
timestamp 1649977179
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1649977179
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1649977179
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_505
timestamp 1649977179
transform 1 0 47564 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_513
timestamp 1649977179
transform 1 0 48300 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_535
timestamp 1649977179
transform 1 0 50324 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_547
timestamp 1649977179
transform 1 0 51428 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1649977179
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1649977179
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1649977179
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_585
timestamp 1649977179
transform 1 0 54924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_597
timestamp 1649977179
transform 1 0 56028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_609
timestamp 1649977179
transform 1 0 57132 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1649977179
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_617
timestamp 1649977179
transform 1 0 57868 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_629
timestamp 1649977179
transform 1 0 58972 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_641
timestamp 1649977179
transform 1 0 60076 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_653
timestamp 1649977179
transform 1 0 61180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_665
timestamp 1649977179
transform 1 0 62284 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_671
timestamp 1649977179
transform 1 0 62836 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_673
timestamp 1649977179
transform 1 0 63020 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_685
timestamp 1649977179
transform 1 0 64124 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_697
timestamp 1649977179
transform 1 0 65228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_709
timestamp 1649977179
transform 1 0 66332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_721
timestamp 1649977179
transform 1 0 67436 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_727
timestamp 1649977179
transform 1 0 67988 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_729
timestamp 1649977179
transform 1 0 68172 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_102_3
timestamp 1649977179
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_15
timestamp 1649977179
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1649977179
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1649977179
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1649977179
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1649977179
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_65
timestamp 1649977179
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1649977179
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1649977179
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_85
timestamp 1649977179
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_97
timestamp 1649977179
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_109
timestamp 1649977179
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_121
timestamp 1649977179
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1649977179
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1649977179
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_141
timestamp 1649977179
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_153
timestamp 1649977179
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_165
timestamp 1649977179
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_177
timestamp 1649977179
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_189
timestamp 1649977179
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1649977179
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_197
timestamp 1649977179
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_209
timestamp 1649977179
transform 1 0 20332 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_221
timestamp 1649977179
transform 1 0 21436 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_233
timestamp 1649977179
transform 1 0 22540 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_245
timestamp 1649977179
transform 1 0 23644 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_251
timestamp 1649977179
transform 1 0 24196 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_253
timestamp 1649977179
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_265
timestamp 1649977179
transform 1 0 25484 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_277
timestamp 1649977179
transform 1 0 26588 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_289
timestamp 1649977179
transform 1 0 27692 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_301
timestamp 1649977179
transform 1 0 28796 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_307
timestamp 1649977179
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_309
timestamp 1649977179
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_321
timestamp 1649977179
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_333
timestamp 1649977179
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_345
timestamp 1649977179
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_357
timestamp 1649977179
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_363
timestamp 1649977179
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_365
timestamp 1649977179
transform 1 0 34684 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_377
timestamp 1649977179
transform 1 0 35788 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_389
timestamp 1649977179
transform 1 0 36892 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_401
timestamp 1649977179
transform 1 0 37996 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_413
timestamp 1649977179
transform 1 0 39100 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_419
timestamp 1649977179
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_421
timestamp 1649977179
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_433
timestamp 1649977179
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_445
timestamp 1649977179
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_457
timestamp 1649977179
transform 1 0 43148 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_469
timestamp 1649977179
transform 1 0 44252 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_475
timestamp 1649977179
transform 1 0 44804 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_477
timestamp 1649977179
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_489
timestamp 1649977179
transform 1 0 46092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_501
timestamp 1649977179
transform 1 0 47196 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_513
timestamp 1649977179
transform 1 0 48300 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_518
timestamp 1649977179
transform 1 0 48760 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_530
timestamp 1649977179
transform 1 0 49864 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_533
timestamp 1649977179
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_545
timestamp 1649977179
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_557
timestamp 1649977179
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_569
timestamp 1649977179
transform 1 0 53452 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_581
timestamp 1649977179
transform 1 0 54556 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_587
timestamp 1649977179
transform 1 0 55108 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_589
timestamp 1649977179
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_601
timestamp 1649977179
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_613
timestamp 1649977179
transform 1 0 57500 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_625
timestamp 1649977179
transform 1 0 58604 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_637
timestamp 1649977179
transform 1 0 59708 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_643
timestamp 1649977179
transform 1 0 60260 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_645
timestamp 1649977179
transform 1 0 60444 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_657
timestamp 1649977179
transform 1 0 61548 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_669
timestamp 1649977179
transform 1 0 62652 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_681
timestamp 1649977179
transform 1 0 63756 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_693
timestamp 1649977179
transform 1 0 64860 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_699
timestamp 1649977179
transform 1 0 65412 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_701
timestamp 1649977179
transform 1 0 65596 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_713
timestamp 1649977179
transform 1 0 66700 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_725
timestamp 1649977179
transform 1 0 67804 0 1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1649977179
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1649977179
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_27
timestamp 1649977179
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_39
timestamp 1649977179
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_51
timestamp 1649977179
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1649977179
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1649977179
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_69
timestamp 1649977179
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_81
timestamp 1649977179
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_93
timestamp 1649977179
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1649977179
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1649977179
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_113
timestamp 1649977179
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_125
timestamp 1649977179
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_137
timestamp 1649977179
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_149
timestamp 1649977179
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_161
timestamp 1649977179
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_167
timestamp 1649977179
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_169
timestamp 1649977179
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_181
timestamp 1649977179
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_193
timestamp 1649977179
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_205
timestamp 1649977179
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_217
timestamp 1649977179
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_223
timestamp 1649977179
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_225
timestamp 1649977179
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_237
timestamp 1649977179
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_249
timestamp 1649977179
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_261
timestamp 1649977179
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_273
timestamp 1649977179
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_279
timestamp 1649977179
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_103_281
timestamp 1649977179
transform 1 0 26956 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_285
timestamp 1649977179
transform 1 0 27324 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_297
timestamp 1649977179
transform 1 0 28428 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_309
timestamp 1649977179
transform 1 0 29532 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_321
timestamp 1649977179
transform 1 0 30636 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_333
timestamp 1649977179
transform 1 0 31740 0 -1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_103_337
timestamp 1649977179
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_349
timestamp 1649977179
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_361
timestamp 1649977179
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_373
timestamp 1649977179
transform 1 0 35420 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_385
timestamp 1649977179
transform 1 0 36524 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_391
timestamp 1649977179
transform 1 0 37076 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_393
timestamp 1649977179
transform 1 0 37260 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_405
timestamp 1649977179
transform 1 0 38364 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_417
timestamp 1649977179
transform 1 0 39468 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_429
timestamp 1649977179
transform 1 0 40572 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_441
timestamp 1649977179
transform 1 0 41676 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_447
timestamp 1649977179
transform 1 0 42228 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_449
timestamp 1649977179
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_461
timestamp 1649977179
transform 1 0 43516 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_473
timestamp 1649977179
transform 1 0 44620 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_485
timestamp 1649977179
transform 1 0 45724 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_497
timestamp 1649977179
transform 1 0 46828 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_503
timestamp 1649977179
transform 1 0 47380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_505
timestamp 1649977179
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_517
timestamp 1649977179
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_529
timestamp 1649977179
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_541
timestamp 1649977179
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_553
timestamp 1649977179
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_559
timestamp 1649977179
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_561
timestamp 1649977179
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_573
timestamp 1649977179
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_585
timestamp 1649977179
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_597
timestamp 1649977179
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_609
timestamp 1649977179
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_615
timestamp 1649977179
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_617
timestamp 1649977179
transform 1 0 57868 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_629
timestamp 1649977179
transform 1 0 58972 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_641
timestamp 1649977179
transform 1 0 60076 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_653
timestamp 1649977179
transform 1 0 61180 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_665
timestamp 1649977179
transform 1 0 62284 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_671
timestamp 1649977179
transform 1 0 62836 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_673
timestamp 1649977179
transform 1 0 63020 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_685
timestamp 1649977179
transform 1 0 64124 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_697
timestamp 1649977179
transform 1 0 65228 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_709
timestamp 1649977179
transform 1 0 66332 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_721
timestamp 1649977179
transform 1 0 67436 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_727
timestamp 1649977179
transform 1 0 67988 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_729
timestamp 1649977179
transform 1 0 68172 0 -1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_104_3
timestamp 1649977179
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_15
timestamp 1649977179
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1649977179
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1649977179
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1649977179
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1649977179
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_65
timestamp 1649977179
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1649977179
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1649977179
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_85
timestamp 1649977179
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_97
timestamp 1649977179
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_109
timestamp 1649977179
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_121
timestamp 1649977179
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1649977179
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1649977179
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_141
timestamp 1649977179
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_153
timestamp 1649977179
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_165
timestamp 1649977179
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_177
timestamp 1649977179
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_189
timestamp 1649977179
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_195
timestamp 1649977179
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_197
timestamp 1649977179
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_209
timestamp 1649977179
transform 1 0 20332 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_221
timestamp 1649977179
transform 1 0 21436 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_233
timestamp 1649977179
transform 1 0 22540 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_245
timestamp 1649977179
transform 1 0 23644 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_251
timestamp 1649977179
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_253
timestamp 1649977179
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_265
timestamp 1649977179
transform 1 0 25484 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_271
timestamp 1649977179
transform 1 0 26036 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_275
timestamp 1649977179
transform 1 0 26404 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_104_300
timestamp 1649977179
transform 1 0 28704 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_104_309
timestamp 1649977179
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_321
timestamp 1649977179
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_333
timestamp 1649977179
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_345
timestamp 1649977179
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_357
timestamp 1649977179
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_363
timestamp 1649977179
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_365
timestamp 1649977179
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_377
timestamp 1649977179
transform 1 0 35788 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_389
timestamp 1649977179
transform 1 0 36892 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_401
timestamp 1649977179
transform 1 0 37996 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_413
timestamp 1649977179
transform 1 0 39100 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_419
timestamp 1649977179
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_421
timestamp 1649977179
transform 1 0 39836 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_433
timestamp 1649977179
transform 1 0 40940 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_445
timestamp 1649977179
transform 1 0 42044 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_457
timestamp 1649977179
transform 1 0 43148 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_469
timestamp 1649977179
transform 1 0 44252 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_475
timestamp 1649977179
transform 1 0 44804 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_477
timestamp 1649977179
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_489
timestamp 1649977179
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_501
timestamp 1649977179
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_513
timestamp 1649977179
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_525
timestamp 1649977179
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_531
timestamp 1649977179
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_533
timestamp 1649977179
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_545
timestamp 1649977179
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_557
timestamp 1649977179
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_569
timestamp 1649977179
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_581
timestamp 1649977179
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_587
timestamp 1649977179
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_589
timestamp 1649977179
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_601
timestamp 1649977179
transform 1 0 56396 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_613
timestamp 1649977179
transform 1 0 57500 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_625
timestamp 1649977179
transform 1 0 58604 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_637
timestamp 1649977179
transform 1 0 59708 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_643
timestamp 1649977179
transform 1 0 60260 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_645
timestamp 1649977179
transform 1 0 60444 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_657
timestamp 1649977179
transform 1 0 61548 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_669
timestamp 1649977179
transform 1 0 62652 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_681
timestamp 1649977179
transform 1 0 63756 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_693
timestamp 1649977179
transform 1 0 64860 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_699
timestamp 1649977179
transform 1 0 65412 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_701
timestamp 1649977179
transform 1 0 65596 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_713
timestamp 1649977179
transform 1 0 66700 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_725
timestamp 1649977179
transform 1 0 67804 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_105_3
timestamp 1649977179
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_15
timestamp 1649977179
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_27
timestamp 1649977179
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_39
timestamp 1649977179
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1649977179
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1649977179
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1649977179
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_69
timestamp 1649977179
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_81
timestamp 1649977179
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_93
timestamp 1649977179
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1649977179
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1649977179
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_113
timestamp 1649977179
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_125
timestamp 1649977179
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_137
timestamp 1649977179
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_149
timestamp 1649977179
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1649977179
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1649977179
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_169
timestamp 1649977179
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_181
timestamp 1649977179
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_193
timestamp 1649977179
transform 1 0 18860 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_205
timestamp 1649977179
transform 1 0 19964 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_217
timestamp 1649977179
transform 1 0 21068 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_223
timestamp 1649977179
transform 1 0 21620 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_225
timestamp 1649977179
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_237
timestamp 1649977179
transform 1 0 22908 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_249
timestamp 1649977179
transform 1 0 24012 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_261
timestamp 1649977179
transform 1 0 25116 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_276
timestamp 1649977179
transform 1 0 26496 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_105_302
timestamp 1649977179
transform 1 0 28888 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_314
timestamp 1649977179
transform 1 0 29992 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_326
timestamp 1649977179
transform 1 0 31096 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_334
timestamp 1649977179
transform 1 0 31832 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_337
timestamp 1649977179
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_349
timestamp 1649977179
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_361
timestamp 1649977179
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_373
timestamp 1649977179
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_385
timestamp 1649977179
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_391
timestamp 1649977179
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_393
timestamp 1649977179
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_405
timestamp 1649977179
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_417
timestamp 1649977179
transform 1 0 39468 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_429
timestamp 1649977179
transform 1 0 40572 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_441
timestamp 1649977179
transform 1 0 41676 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_447
timestamp 1649977179
transform 1 0 42228 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_449
timestamp 1649977179
transform 1 0 42412 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_461
timestamp 1649977179
transform 1 0 43516 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_473
timestamp 1649977179
transform 1 0 44620 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_485
timestamp 1649977179
transform 1 0 45724 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_497
timestamp 1649977179
transform 1 0 46828 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_503
timestamp 1649977179
transform 1 0 47380 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_508
timestamp 1649977179
transform 1 0 47840 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_520
timestamp 1649977179
transform 1 0 48944 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_532
timestamp 1649977179
transform 1 0 50048 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_544
timestamp 1649977179
transform 1 0 51152 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_556
timestamp 1649977179
transform 1 0 52256 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_105_561
timestamp 1649977179
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_573
timestamp 1649977179
transform 1 0 53820 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_585
timestamp 1649977179
transform 1 0 54924 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_597
timestamp 1649977179
transform 1 0 56028 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_609
timestamp 1649977179
transform 1 0 57132 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_615
timestamp 1649977179
transform 1 0 57684 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_617
timestamp 1649977179
transform 1 0 57868 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_629
timestamp 1649977179
transform 1 0 58972 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_641
timestamp 1649977179
transform 1 0 60076 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_653
timestamp 1649977179
transform 1 0 61180 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_665
timestamp 1649977179
transform 1 0 62284 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_671
timestamp 1649977179
transform 1 0 62836 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_673
timestamp 1649977179
transform 1 0 63020 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_685
timestamp 1649977179
transform 1 0 64124 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_697
timestamp 1649977179
transform 1 0 65228 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_709
timestamp 1649977179
transform 1 0 66332 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_721
timestamp 1649977179
transform 1 0 67436 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_727
timestamp 1649977179
transform 1 0 67988 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_729
timestamp 1649977179
transform 1 0 68172 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1649977179
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1649977179
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1649977179
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1649977179
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1649977179
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1649977179
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_65
timestamp 1649977179
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1649977179
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1649977179
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_85
timestamp 1649977179
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_97
timestamp 1649977179
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_109
timestamp 1649977179
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_121
timestamp 1649977179
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_133
timestamp 1649977179
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1649977179
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_141
timestamp 1649977179
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_153
timestamp 1649977179
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_165
timestamp 1649977179
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_177
timestamp 1649977179
transform 1 0 17388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_189
timestamp 1649977179
transform 1 0 18492 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_195
timestamp 1649977179
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_197
timestamp 1649977179
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_209
timestamp 1649977179
transform 1 0 20332 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_221
timestamp 1649977179
transform 1 0 21436 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_233
timestamp 1649977179
transform 1 0 22540 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_241
timestamp 1649977179
transform 1 0 23276 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_106_246
timestamp 1649977179
transform 1 0 23736 0 1 59840
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_106_253
timestamp 1649977179
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_265
timestamp 1649977179
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_277
timestamp 1649977179
transform 1 0 26588 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_282
timestamp 1649977179
transform 1 0 27048 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_294
timestamp 1649977179
transform 1 0 28152 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_306
timestamp 1649977179
transform 1 0 29256 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_309
timestamp 1649977179
transform 1 0 29532 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_321
timestamp 1649977179
transform 1 0 30636 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_333
timestamp 1649977179
transform 1 0 31740 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_345
timestamp 1649977179
transform 1 0 32844 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_357
timestamp 1649977179
transform 1 0 33948 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_363
timestamp 1649977179
transform 1 0 34500 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_365
timestamp 1649977179
transform 1 0 34684 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_377
timestamp 1649977179
transform 1 0 35788 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_389
timestamp 1649977179
transform 1 0 36892 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_401
timestamp 1649977179
transform 1 0 37996 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_413
timestamp 1649977179
transform 1 0 39100 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_419
timestamp 1649977179
transform 1 0 39652 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_421
timestamp 1649977179
transform 1 0 39836 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_433
timestamp 1649977179
transform 1 0 40940 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_445
timestamp 1649977179
transform 1 0 42044 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_457
timestamp 1649977179
transform 1 0 43148 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_469
timestamp 1649977179
transform 1 0 44252 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_475
timestamp 1649977179
transform 1 0 44804 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_477
timestamp 1649977179
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_489
timestamp 1649977179
transform 1 0 46092 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_496
timestamp 1649977179
transform 1 0 46736 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_521
timestamp 1649977179
transform 1 0 49036 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_106_529
timestamp 1649977179
transform 1 0 49772 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_533
timestamp 1649977179
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_545
timestamp 1649977179
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_557
timestamp 1649977179
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_569
timestamp 1649977179
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_581
timestamp 1649977179
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_587
timestamp 1649977179
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_589
timestamp 1649977179
transform 1 0 55292 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_601
timestamp 1649977179
transform 1 0 56396 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_613
timestamp 1649977179
transform 1 0 57500 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_625
timestamp 1649977179
transform 1 0 58604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_637
timestamp 1649977179
transform 1 0 59708 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_643
timestamp 1649977179
transform 1 0 60260 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_645
timestamp 1649977179
transform 1 0 60444 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_657
timestamp 1649977179
transform 1 0 61548 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_669
timestamp 1649977179
transform 1 0 62652 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_681
timestamp 1649977179
transform 1 0 63756 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_693
timestamp 1649977179
transform 1 0 64860 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_699
timestamp 1649977179
transform 1 0 65412 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_701
timestamp 1649977179
transform 1 0 65596 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_713
timestamp 1649977179
transform 1 0 66700 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_725
timestamp 1649977179
transform 1 0 67804 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_107_13
timestamp 1649977179
transform 1 0 2300 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_25
timestamp 1649977179
transform 1 0 3404 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_37
timestamp 1649977179
transform 1 0 4508 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_49
timestamp 1649977179
transform 1 0 5612 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1649977179
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1649977179
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_69
timestamp 1649977179
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_81
timestamp 1649977179
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_93
timestamp 1649977179
transform 1 0 9660 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_105
timestamp 1649977179
transform 1 0 10764 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_111
timestamp 1649977179
transform 1 0 11316 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_113
timestamp 1649977179
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_125
timestamp 1649977179
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_137
timestamp 1649977179
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_149
timestamp 1649977179
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_161
timestamp 1649977179
transform 1 0 15916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_167
timestamp 1649977179
transform 1 0 16468 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_169
timestamp 1649977179
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_181
timestamp 1649977179
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_193
timestamp 1649977179
transform 1 0 18860 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_205
timestamp 1649977179
transform 1 0 19964 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_217
timestamp 1649977179
transform 1 0 21068 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_223
timestamp 1649977179
transform 1 0 21620 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_225
timestamp 1649977179
transform 1 0 21804 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_237
timestamp 1649977179
transform 1 0 22908 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_259
timestamp 1649977179
transform 1 0 24932 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_271
timestamp 1649977179
transform 1 0 26036 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_279
timestamp 1649977179
transform 1 0 26772 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_281
timestamp 1649977179
transform 1 0 26956 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_293
timestamp 1649977179
transform 1 0 28060 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_305
timestamp 1649977179
transform 1 0 29164 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_317
timestamp 1649977179
transform 1 0 30268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_329
timestamp 1649977179
transform 1 0 31372 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_335
timestamp 1649977179
transform 1 0 31924 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_337
timestamp 1649977179
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_349
timestamp 1649977179
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_361
timestamp 1649977179
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_373
timestamp 1649977179
transform 1 0 35420 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_385
timestamp 1649977179
transform 1 0 36524 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_391
timestamp 1649977179
transform 1 0 37076 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_393
timestamp 1649977179
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_405
timestamp 1649977179
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_417
timestamp 1649977179
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_429
timestamp 1649977179
transform 1 0 40572 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_441
timestamp 1649977179
transform 1 0 41676 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_447
timestamp 1649977179
transform 1 0 42228 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_449
timestamp 1649977179
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_461
timestamp 1649977179
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_473
timestamp 1649977179
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_485
timestamp 1649977179
transform 1 0 45724 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_497
timestamp 1649977179
transform 1 0 46828 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_503
timestamp 1649977179
transform 1 0 47380 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_505
timestamp 1649977179
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_517
timestamp 1649977179
transform 1 0 48668 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_529
timestamp 1649977179
transform 1 0 49772 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_541
timestamp 1649977179
transform 1 0 50876 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_553
timestamp 1649977179
transform 1 0 51980 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_559
timestamp 1649977179
transform 1 0 52532 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_561
timestamp 1649977179
transform 1 0 52716 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_573
timestamp 1649977179
transform 1 0 53820 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_585
timestamp 1649977179
transform 1 0 54924 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_597
timestamp 1649977179
transform 1 0 56028 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_609
timestamp 1649977179
transform 1 0 57132 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_615
timestamp 1649977179
transform 1 0 57684 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_617
timestamp 1649977179
transform 1 0 57868 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_629
timestamp 1649977179
transform 1 0 58972 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_641
timestamp 1649977179
transform 1 0 60076 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_653
timestamp 1649977179
transform 1 0 61180 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_665
timestamp 1649977179
transform 1 0 62284 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_671
timestamp 1649977179
transform 1 0 62836 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_673
timestamp 1649977179
transform 1 0 63020 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_685
timestamp 1649977179
transform 1 0 64124 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_697
timestamp 1649977179
transform 1 0 65228 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_709
timestamp 1649977179
transform 1 0 66332 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_721
timestamp 1649977179
transform 1 0 67436 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_727
timestamp 1649977179
transform 1 0 67988 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_729
timestamp 1649977179
transform 1 0 68172 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1649977179
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1649977179
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1649977179
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1649977179
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_41
timestamp 1649977179
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_53
timestamp 1649977179
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_65
timestamp 1649977179
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1649977179
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1649977179
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_85
timestamp 1649977179
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_97
timestamp 1649977179
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_109
timestamp 1649977179
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_121
timestamp 1649977179
transform 1 0 12236 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_133
timestamp 1649977179
transform 1 0 13340 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_139
timestamp 1649977179
transform 1 0 13892 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_141
timestamp 1649977179
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_153
timestamp 1649977179
transform 1 0 15180 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_165
timestamp 1649977179
transform 1 0 16284 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_177
timestamp 1649977179
transform 1 0 17388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_189
timestamp 1649977179
transform 1 0 18492 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_195
timestamp 1649977179
transform 1 0 19044 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_197
timestamp 1649977179
transform 1 0 19228 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_209
timestamp 1649977179
transform 1 0 20332 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_221
timestamp 1649977179
transform 1 0 21436 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_108_233
timestamp 1649977179
transform 1 0 22540 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_237
timestamp 1649977179
transform 1 0 22908 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_241
timestamp 1649977179
transform 1 0 23276 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_108_249
timestamp 1649977179
transform 1 0 24012 0 1 60928
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_108_253
timestamp 1649977179
transform 1 0 24380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_265
timestamp 1649977179
transform 1 0 25484 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_277
timestamp 1649977179
transform 1 0 26588 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_289
timestamp 1649977179
transform 1 0 27692 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_301
timestamp 1649977179
transform 1 0 28796 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_307
timestamp 1649977179
transform 1 0 29348 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_309
timestamp 1649977179
transform 1 0 29532 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_321
timestamp 1649977179
transform 1 0 30636 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_333
timestamp 1649977179
transform 1 0 31740 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_345
timestamp 1649977179
transform 1 0 32844 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_357
timestamp 1649977179
transform 1 0 33948 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_363
timestamp 1649977179
transform 1 0 34500 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_365
timestamp 1649977179
transform 1 0 34684 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_377
timestamp 1649977179
transform 1 0 35788 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_389
timestamp 1649977179
transform 1 0 36892 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_401
timestamp 1649977179
transform 1 0 37996 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_413
timestamp 1649977179
transform 1 0 39100 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_419
timestamp 1649977179
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_421
timestamp 1649977179
transform 1 0 39836 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_433
timestamp 1649977179
transform 1 0 40940 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_445
timestamp 1649977179
transform 1 0 42044 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_457
timestamp 1649977179
transform 1 0 43148 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_469
timestamp 1649977179
transform 1 0 44252 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_475
timestamp 1649977179
transform 1 0 44804 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_477
timestamp 1649977179
transform 1 0 44988 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_489
timestamp 1649977179
transform 1 0 46092 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_501
timestamp 1649977179
transform 1 0 47196 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_513
timestamp 1649977179
transform 1 0 48300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_525
timestamp 1649977179
transform 1 0 49404 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1649977179
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_533
timestamp 1649977179
transform 1 0 50140 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_545
timestamp 1649977179
transform 1 0 51244 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_557
timestamp 1649977179
transform 1 0 52348 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_569
timestamp 1649977179
transform 1 0 53452 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_577
timestamp 1649977179
transform 1 0 54188 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_108_582
timestamp 1649977179
transform 1 0 54648 0 1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_108_589
timestamp 1649977179
transform 1 0 55292 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_601
timestamp 1649977179
transform 1 0 56396 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_613
timestamp 1649977179
transform 1 0 57500 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_625
timestamp 1649977179
transform 1 0 58604 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_637
timestamp 1649977179
transform 1 0 59708 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_643
timestamp 1649977179
transform 1 0 60260 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_645
timestamp 1649977179
transform 1 0 60444 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_657
timestamp 1649977179
transform 1 0 61548 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_669
timestamp 1649977179
transform 1 0 62652 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_681
timestamp 1649977179
transform 1 0 63756 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_693
timestamp 1649977179
transform 1 0 64860 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_699
timestamp 1649977179
transform 1 0 65412 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_701
timestamp 1649977179
transform 1 0 65596 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_713
timestamp 1649977179
transform 1 0 66700 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_725
timestamp 1649977179
transform 1 0 67804 0 1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_109_3
timestamp 1649977179
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_15
timestamp 1649977179
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_27
timestamp 1649977179
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_39
timestamp 1649977179
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1649977179
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1649977179
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_57
timestamp 1649977179
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_69
timestamp 1649977179
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_81
timestamp 1649977179
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_93
timestamp 1649977179
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_105
timestamp 1649977179
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_111
timestamp 1649977179
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_113
timestamp 1649977179
transform 1 0 11500 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_125
timestamp 1649977179
transform 1 0 12604 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_137
timestamp 1649977179
transform 1 0 13708 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_149
timestamp 1649977179
transform 1 0 14812 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_161
timestamp 1649977179
transform 1 0 15916 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_167
timestamp 1649977179
transform 1 0 16468 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_169
timestamp 1649977179
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_181
timestamp 1649977179
transform 1 0 17756 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_193
timestamp 1649977179
transform 1 0 18860 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_205
timestamp 1649977179
transform 1 0 19964 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_217
timestamp 1649977179
transform 1 0 21068 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_223
timestamp 1649977179
transform 1 0 21620 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_225
timestamp 1649977179
transform 1 0 21804 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_237
timestamp 1649977179
transform 1 0 22908 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_249
timestamp 1649977179
transform 1 0 24012 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_261
timestamp 1649977179
transform 1 0 25116 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_273
timestamp 1649977179
transform 1 0 26220 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_279
timestamp 1649977179
transform 1 0 26772 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_281
timestamp 1649977179
transform 1 0 26956 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_293
timestamp 1649977179
transform 1 0 28060 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_305
timestamp 1649977179
transform 1 0 29164 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_317
timestamp 1649977179
transform 1 0 30268 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_329
timestamp 1649977179
transform 1 0 31372 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_335
timestamp 1649977179
transform 1 0 31924 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_337
timestamp 1649977179
transform 1 0 32108 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_349
timestamp 1649977179
transform 1 0 33212 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_361
timestamp 1649977179
transform 1 0 34316 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_373
timestamp 1649977179
transform 1 0 35420 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_385
timestamp 1649977179
transform 1 0 36524 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_391
timestamp 1649977179
transform 1 0 37076 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_393
timestamp 1649977179
transform 1 0 37260 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_405
timestamp 1649977179
transform 1 0 38364 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_417
timestamp 1649977179
transform 1 0 39468 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_429
timestamp 1649977179
transform 1 0 40572 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_441
timestamp 1649977179
transform 1 0 41676 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_447
timestamp 1649977179
transform 1 0 42228 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_449
timestamp 1649977179
transform 1 0 42412 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_461
timestamp 1649977179
transform 1 0 43516 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_473
timestamp 1649977179
transform 1 0 44620 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_485
timestamp 1649977179
transform 1 0 45724 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_109_493
timestamp 1649977179
transform 1 0 46460 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_109_497
timestamp 1649977179
transform 1 0 46828 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_503
timestamp 1649977179
transform 1 0 47380 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_505
timestamp 1649977179
transform 1 0 47564 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_517
timestamp 1649977179
transform 1 0 48668 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_529
timestamp 1649977179
transform 1 0 49772 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_541
timestamp 1649977179
transform 1 0 50876 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_553
timestamp 1649977179
transform 1 0 51980 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_559
timestamp 1649977179
transform 1 0 52532 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_561
timestamp 1649977179
transform 1 0 52716 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_573
timestamp 1649977179
transform 1 0 53820 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_579
timestamp 1649977179
transform 1 0 54372 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_601
timestamp 1649977179
transform 1 0 56396 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_109_613
timestamp 1649977179
transform 1 0 57500 0 -1 62016
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_109_617
timestamp 1649977179
transform 1 0 57868 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_629
timestamp 1649977179
transform 1 0 58972 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_641
timestamp 1649977179
transform 1 0 60076 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_653
timestamp 1649977179
transform 1 0 61180 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_665
timestamp 1649977179
transform 1 0 62284 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_671
timestamp 1649977179
transform 1 0 62836 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_673
timestamp 1649977179
transform 1 0 63020 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_685
timestamp 1649977179
transform 1 0 64124 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_692
timestamp 1649977179
transform 1 0 64768 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_109_717
timestamp 1649977179
transform 1 0 67068 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_109_725
timestamp 1649977179
transform 1 0 67804 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_109_729
timestamp 1649977179
transform 1 0 68172 0 -1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_110_3
timestamp 1649977179
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_15
timestamp 1649977179
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1649977179
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1649977179
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_41
timestamp 1649977179
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_53
timestamp 1649977179
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_65
timestamp 1649977179
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1649977179
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1649977179
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_85
timestamp 1649977179
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_97
timestamp 1649977179
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_109
timestamp 1649977179
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_121
timestamp 1649977179
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_133
timestamp 1649977179
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_139
timestamp 1649977179
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_141
timestamp 1649977179
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_153
timestamp 1649977179
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_165
timestamp 1649977179
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_177
timestamp 1649977179
transform 1 0 17388 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_189
timestamp 1649977179
transform 1 0 18492 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_195
timestamp 1649977179
transform 1 0 19044 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_197
timestamp 1649977179
transform 1 0 19228 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_209
timestamp 1649977179
transform 1 0 20332 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_221
timestamp 1649977179
transform 1 0 21436 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_233
timestamp 1649977179
transform 1 0 22540 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_245
timestamp 1649977179
transform 1 0 23644 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_251
timestamp 1649977179
transform 1 0 24196 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_253
timestamp 1649977179
transform 1 0 24380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_265
timestamp 1649977179
transform 1 0 25484 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_277
timestamp 1649977179
transform 1 0 26588 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_289
timestamp 1649977179
transform 1 0 27692 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_301
timestamp 1649977179
transform 1 0 28796 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_307
timestamp 1649977179
transform 1 0 29348 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_309
timestamp 1649977179
transform 1 0 29532 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_321
timestamp 1649977179
transform 1 0 30636 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_333
timestamp 1649977179
transform 1 0 31740 0 1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_110_342
timestamp 1649977179
transform 1 0 32568 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_354
timestamp 1649977179
transform 1 0 33672 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_110_362
timestamp 1649977179
transform 1 0 34408 0 1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_110_365
timestamp 1649977179
transform 1 0 34684 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_377
timestamp 1649977179
transform 1 0 35788 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_389
timestamp 1649977179
transform 1 0 36892 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_401
timestamp 1649977179
transform 1 0 37996 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_413
timestamp 1649977179
transform 1 0 39100 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_419
timestamp 1649977179
transform 1 0 39652 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_421
timestamp 1649977179
transform 1 0 39836 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_433
timestamp 1649977179
transform 1 0 40940 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_445
timestamp 1649977179
transform 1 0 42044 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_457
timestamp 1649977179
transform 1 0 43148 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_469
timestamp 1649977179
transform 1 0 44252 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_475
timestamp 1649977179
transform 1 0 44804 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_477
timestamp 1649977179
transform 1 0 44988 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_489
timestamp 1649977179
transform 1 0 46092 0 1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_110_514
timestamp 1649977179
transform 1 0 48392 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_526
timestamp 1649977179
transform 1 0 49496 0 1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_110_536
timestamp 1649977179
transform 1 0 50416 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_548
timestamp 1649977179
transform 1 0 51520 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_560
timestamp 1649977179
transform 1 0 52624 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_572
timestamp 1649977179
transform 1 0 53728 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_110_583
timestamp 1649977179
transform 1 0 54740 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_587
timestamp 1649977179
transform 1 0 55108 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_589
timestamp 1649977179
transform 1 0 55292 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_601
timestamp 1649977179
transform 1 0 56396 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_613
timestamp 1649977179
transform 1 0 57500 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_625
timestamp 1649977179
transform 1 0 58604 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_637
timestamp 1649977179
transform 1 0 59708 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_643
timestamp 1649977179
transform 1 0 60260 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_645
timestamp 1649977179
transform 1 0 60444 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_657
timestamp 1649977179
transform 1 0 61548 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_669
timestamp 1649977179
transform 1 0 62652 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_681
timestamp 1649977179
transform 1 0 63756 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_696
timestamp 1649977179
transform 1 0 65136 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_110_722
timestamp 1649977179
transform 1 0 67528 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_110_730
timestamp 1649977179
transform 1 0 68264 0 1 62016
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1649977179
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1649977179
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_27
timestamp 1649977179
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_39
timestamp 1649977179
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1649977179
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1649977179
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_57
timestamp 1649977179
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_69
timestamp 1649977179
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_81
timestamp 1649977179
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_93
timestamp 1649977179
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_105
timestamp 1649977179
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_111
timestamp 1649977179
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_113
timestamp 1649977179
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_125
timestamp 1649977179
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_137
timestamp 1649977179
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_149
timestamp 1649977179
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_161
timestamp 1649977179
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_167
timestamp 1649977179
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_169
timestamp 1649977179
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_181
timestamp 1649977179
transform 1 0 17756 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_193
timestamp 1649977179
transform 1 0 18860 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_205
timestamp 1649977179
transform 1 0 19964 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_217
timestamp 1649977179
transform 1 0 21068 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_223
timestamp 1649977179
transform 1 0 21620 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_225
timestamp 1649977179
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_237
timestamp 1649977179
transform 1 0 22908 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_249
timestamp 1649977179
transform 1 0 24012 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_261
timestamp 1649977179
transform 1 0 25116 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_273
timestamp 1649977179
transform 1 0 26220 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_279
timestamp 1649977179
transform 1 0 26772 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_281
timestamp 1649977179
transform 1 0 26956 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_293
timestamp 1649977179
transform 1 0 28060 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_305
timestamp 1649977179
transform 1 0 29164 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_317
timestamp 1649977179
transform 1 0 30268 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_332
timestamp 1649977179
transform 1 0 31648 0 -1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_111_358
timestamp 1649977179
transform 1 0 34040 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_370
timestamp 1649977179
transform 1 0 35144 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_382
timestamp 1649977179
transform 1 0 36248 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_111_390
timestamp 1649977179
transform 1 0 36984 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_111_393
timestamp 1649977179
transform 1 0 37260 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_405
timestamp 1649977179
transform 1 0 38364 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_417
timestamp 1649977179
transform 1 0 39468 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_429
timestamp 1649977179
transform 1 0 40572 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_441
timestamp 1649977179
transform 1 0 41676 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_447
timestamp 1649977179
transform 1 0 42228 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_449
timestamp 1649977179
transform 1 0 42412 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_461
timestamp 1649977179
transform 1 0 43516 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_473
timestamp 1649977179
transform 1 0 44620 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_485
timestamp 1649977179
transform 1 0 45724 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_493
timestamp 1649977179
transform 1 0 46460 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_111_497
timestamp 1649977179
transform 1 0 46828 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_503
timestamp 1649977179
transform 1 0 47380 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_505
timestamp 1649977179
transform 1 0 47564 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_517
timestamp 1649977179
transform 1 0 48668 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_111_524
timestamp 1649977179
transform 1 0 49312 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_111_549
timestamp 1649977179
transform 1 0 51612 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_111_557
timestamp 1649977179
transform 1 0 52348 0 -1 63104
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_111_561
timestamp 1649977179
transform 1 0 52716 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_573
timestamp 1649977179
transform 1 0 53820 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_585
timestamp 1649977179
transform 1 0 54924 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_597
timestamp 1649977179
transform 1 0 56028 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_609
timestamp 1649977179
transform 1 0 57132 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_615
timestamp 1649977179
transform 1 0 57684 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_620
timestamp 1649977179
transform 1 0 58144 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_632
timestamp 1649977179
transform 1 0 59248 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_644
timestamp 1649977179
transform 1 0 60352 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_656
timestamp 1649977179
transform 1 0 61456 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_668
timestamp 1649977179
transform 1 0 62560 0 -1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_111_673
timestamp 1649977179
transform 1 0 63020 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_685
timestamp 1649977179
transform 1 0 64124 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_693
timestamp 1649977179
transform 1 0 64860 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_111_697
timestamp 1649977179
transform 1 0 65228 0 -1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_111_704
timestamp 1649977179
transform 1 0 65872 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_716
timestamp 1649977179
transform 1 0 66976 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_729
timestamp 1649977179
transform 1 0 68172 0 -1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_112_3
timestamp 1649977179
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_15
timestamp 1649977179
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1649977179
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1649977179
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_41
timestamp 1649977179
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_53
timestamp 1649977179
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_65
timestamp 1649977179
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1649977179
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1649977179
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_85
timestamp 1649977179
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_97
timestamp 1649977179
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_109
timestamp 1649977179
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_121
timestamp 1649977179
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_133
timestamp 1649977179
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_139
timestamp 1649977179
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_141
timestamp 1649977179
transform 1 0 14076 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_153
timestamp 1649977179
transform 1 0 15180 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_165
timestamp 1649977179
transform 1 0 16284 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_177
timestamp 1649977179
transform 1 0 17388 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_189
timestamp 1649977179
transform 1 0 18492 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_195
timestamp 1649977179
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_197
timestamp 1649977179
transform 1 0 19228 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_209
timestamp 1649977179
transform 1 0 20332 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_221
timestamp 1649977179
transform 1 0 21436 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_233
timestamp 1649977179
transform 1 0 22540 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_245
timestamp 1649977179
transform 1 0 23644 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_251
timestamp 1649977179
transform 1 0 24196 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_253
timestamp 1649977179
transform 1 0 24380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_265
timestamp 1649977179
transform 1 0 25484 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_277
timestamp 1649977179
transform 1 0 26588 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_289
timestamp 1649977179
transform 1 0 27692 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_301
timestamp 1649977179
transform 1 0 28796 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_307
timestamp 1649977179
transform 1 0 29348 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_309
timestamp 1649977179
transform 1 0 29532 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_112_324
timestamp 1649977179
transform 1 0 30912 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_344
timestamp 1649977179
transform 1 0 32752 0 1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_112_351
timestamp 1649977179
transform 1 0 33396 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_363
timestamp 1649977179
transform 1 0 34500 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_365
timestamp 1649977179
transform 1 0 34684 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_377
timestamp 1649977179
transform 1 0 35788 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_389
timestamp 1649977179
transform 1 0 36892 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_401
timestamp 1649977179
transform 1 0 37996 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_413
timestamp 1649977179
transform 1 0 39100 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_419
timestamp 1649977179
transform 1 0 39652 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_421
timestamp 1649977179
transform 1 0 39836 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_433
timestamp 1649977179
transform 1 0 40940 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_445
timestamp 1649977179
transform 1 0 42044 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_457
timestamp 1649977179
transform 1 0 43148 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_469
timestamp 1649977179
transform 1 0 44252 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_475
timestamp 1649977179
transform 1 0 44804 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_477
timestamp 1649977179
transform 1 0 44988 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_489
timestamp 1649977179
transform 1 0 46092 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_501
timestamp 1649977179
transform 1 0 47196 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_513
timestamp 1649977179
transform 1 0 48300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_525
timestamp 1649977179
transform 1 0 49404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_531
timestamp 1649977179
transform 1 0 49956 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_536
timestamp 1649977179
transform 1 0 50416 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_548
timestamp 1649977179
transform 1 0 51520 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_560
timestamp 1649977179
transform 1 0 52624 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_572
timestamp 1649977179
transform 1 0 53728 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_112_584
timestamp 1649977179
transform 1 0 54832 0 1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_112_589
timestamp 1649977179
transform 1 0 55292 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_601
timestamp 1649977179
transform 1 0 56396 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_613
timestamp 1649977179
transform 1 0 57500 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_635
timestamp 1649977179
transform 1 0 59524 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_112_643
timestamp 1649977179
transform 1 0 60260 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_645
timestamp 1649977179
transform 1 0 60444 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_657
timestamp 1649977179
transform 1 0 61548 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_669
timestamp 1649977179
transform 1 0 62652 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_681
timestamp 1649977179
transform 1 0 63756 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_693
timestamp 1649977179
transform 1 0 64860 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_699
timestamp 1649977179
transform 1 0 65412 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_701
timestamp 1649977179
transform 1 0 65596 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_713
timestamp 1649977179
transform 1 0 66700 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_725
timestamp 1649977179
transform 1 0 67804 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1649977179
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1649977179
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1649977179
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_39
timestamp 1649977179
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1649977179
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1649977179
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_57
timestamp 1649977179
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_69
timestamp 1649977179
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_81
timestamp 1649977179
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_93
timestamp 1649977179
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_105
timestamp 1649977179
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_111
timestamp 1649977179
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_113
timestamp 1649977179
transform 1 0 11500 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_125
timestamp 1649977179
transform 1 0 12604 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_137
timestamp 1649977179
transform 1 0 13708 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_149
timestamp 1649977179
transform 1 0 14812 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_161
timestamp 1649977179
transform 1 0 15916 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_167
timestamp 1649977179
transform 1 0 16468 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_169
timestamp 1649977179
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_181
timestamp 1649977179
transform 1 0 17756 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_193
timestamp 1649977179
transform 1 0 18860 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_205
timestamp 1649977179
transform 1 0 19964 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_217
timestamp 1649977179
transform 1 0 21068 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_223
timestamp 1649977179
transform 1 0 21620 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_225
timestamp 1649977179
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_237
timestamp 1649977179
transform 1 0 22908 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_249
timestamp 1649977179
transform 1 0 24012 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_261
timestamp 1649977179
transform 1 0 25116 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_273
timestamp 1649977179
transform 1 0 26220 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_279
timestamp 1649977179
transform 1 0 26772 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_281
timestamp 1649977179
transform 1 0 26956 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_293
timestamp 1649977179
transform 1 0 28060 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_113_302
timestamp 1649977179
transform 1 0 28888 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_113_327
timestamp 1649977179
transform 1 0 31188 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_113_335
timestamp 1649977179
transform 1 0 31924 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_358
timestamp 1649977179
transform 1 0 34040 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_370
timestamp 1649977179
transform 1 0 35144 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_382
timestamp 1649977179
transform 1 0 36248 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_113_390
timestamp 1649977179
transform 1 0 36984 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_113_393
timestamp 1649977179
transform 1 0 37260 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_405
timestamp 1649977179
transform 1 0 38364 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_417
timestamp 1649977179
transform 1 0 39468 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_429
timestamp 1649977179
transform 1 0 40572 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_441
timestamp 1649977179
transform 1 0 41676 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_447
timestamp 1649977179
transform 1 0 42228 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_449
timestamp 1649977179
transform 1 0 42412 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_461
timestamp 1649977179
transform 1 0 43516 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_473
timestamp 1649977179
transform 1 0 44620 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_485
timestamp 1649977179
transform 1 0 45724 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_497
timestamp 1649977179
transform 1 0 46828 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_503
timestamp 1649977179
transform 1 0 47380 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_505
timestamp 1649977179
transform 1 0 47564 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_517
timestamp 1649977179
transform 1 0 48668 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_529
timestamp 1649977179
transform 1 0 49772 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_541
timestamp 1649977179
transform 1 0 50876 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_553
timestamp 1649977179
transform 1 0 51980 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_559
timestamp 1649977179
transform 1 0 52532 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_561
timestamp 1649977179
transform 1 0 52716 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_573
timestamp 1649977179
transform 1 0 53820 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_585
timestamp 1649977179
transform 1 0 54924 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_591
timestamp 1649977179
transform 1 0 55476 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_595
timestamp 1649977179
transform 1 0 55844 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_607
timestamp 1649977179
transform 1 0 56948 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_113_615
timestamp 1649977179
transform 1 0 57684 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_620
timestamp 1649977179
transform 1 0 58144 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_632
timestamp 1649977179
transform 1 0 59248 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_644
timestamp 1649977179
transform 1 0 60352 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_656
timestamp 1649977179
transform 1 0 61456 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_668
timestamp 1649977179
transform 1 0 62560 0 -1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_113_673
timestamp 1649977179
transform 1 0 63020 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_685
timestamp 1649977179
transform 1 0 64124 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_697
timestamp 1649977179
transform 1 0 65228 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_709
timestamp 1649977179
transform 1 0 66332 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_721
timestamp 1649977179
transform 1 0 67436 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_727
timestamp 1649977179
transform 1 0 67988 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_113_729
timestamp 1649977179
transform 1 0 68172 0 -1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_114_3
timestamp 1649977179
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_15
timestamp 1649977179
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1649977179
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1649977179
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_41
timestamp 1649977179
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_53
timestamp 1649977179
transform 1 0 5980 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_114_61
timestamp 1649977179
transform 1 0 6716 0 1 64192
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_114_67
timestamp 1649977179
transform 1 0 7268 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_114_79
timestamp 1649977179
transform 1 0 8372 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1649977179
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_85
timestamp 1649977179
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_97
timestamp 1649977179
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_109
timestamp 1649977179
transform 1 0 11132 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_121
timestamp 1649977179
transform 1 0 12236 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_133
timestamp 1649977179
transform 1 0 13340 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_139
timestamp 1649977179
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_141
timestamp 1649977179
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_153
timestamp 1649977179
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_165
timestamp 1649977179
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_177
timestamp 1649977179
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_189
timestamp 1649977179
transform 1 0 18492 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_195
timestamp 1649977179
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_197
timestamp 1649977179
transform 1 0 19228 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_209
timestamp 1649977179
transform 1 0 20332 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_221
timestamp 1649977179
transform 1 0 21436 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_233
timestamp 1649977179
transform 1 0 22540 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_245
timestamp 1649977179
transform 1 0 23644 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_251
timestamp 1649977179
transform 1 0 24196 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_253
timestamp 1649977179
transform 1 0 24380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_265
timestamp 1649977179
transform 1 0 25484 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_277
timestamp 1649977179
transform 1 0 26588 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_289
timestamp 1649977179
transform 1 0 27692 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_301
timestamp 1649977179
transform 1 0 28796 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_307
timestamp 1649977179
transform 1 0 29348 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_114_312
timestamp 1649977179
transform 1 0 29808 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_114_317
timestamp 1649977179
transform 1 0 30268 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_114_321
timestamp 1649977179
transform 1 0 30636 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_114_328
timestamp 1649977179
transform 1 0 31280 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_353
timestamp 1649977179
transform 1 0 33580 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_360
timestamp 1649977179
transform 1 0 34224 0 1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_114_365
timestamp 1649977179
transform 1 0 34684 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_377
timestamp 1649977179
transform 1 0 35788 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_389
timestamp 1649977179
transform 1 0 36892 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_401
timestamp 1649977179
transform 1 0 37996 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_413
timestamp 1649977179
transform 1 0 39100 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_419
timestamp 1649977179
transform 1 0 39652 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_421
timestamp 1649977179
transform 1 0 39836 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_433
timestamp 1649977179
transform 1 0 40940 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_445
timestamp 1649977179
transform 1 0 42044 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_451
timestamp 1649977179
transform 1 0 42596 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_455
timestamp 1649977179
transform 1 0 42964 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_467
timestamp 1649977179
transform 1 0 44068 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_114_475
timestamp 1649977179
transform 1 0 44804 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_477
timestamp 1649977179
transform 1 0 44988 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_489
timestamp 1649977179
transform 1 0 46092 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_501
timestamp 1649977179
transform 1 0 47196 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_513
timestamp 1649977179
transform 1 0 48300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_525
timestamp 1649977179
transform 1 0 49404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_531
timestamp 1649977179
transform 1 0 49956 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_533
timestamp 1649977179
transform 1 0 50140 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_545
timestamp 1649977179
transform 1 0 51244 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_557
timestamp 1649977179
transform 1 0 52348 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_569
timestamp 1649977179
transform 1 0 53452 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_581
timestamp 1649977179
transform 1 0 54556 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_587
timestamp 1649977179
transform 1 0 55108 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_114_589
timestamp 1649977179
transform 1 0 55292 0 1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_114_614
timestamp 1649977179
transform 1 0 57592 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_626
timestamp 1649977179
transform 1 0 58696 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_638
timestamp 1649977179
transform 1 0 59800 0 1 64192
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_114_645
timestamp 1649977179
transform 1 0 60444 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_657
timestamp 1649977179
transform 1 0 61548 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_669
timestamp 1649977179
transform 1 0 62652 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_681
timestamp 1649977179
transform 1 0 63756 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_693
timestamp 1649977179
transform 1 0 64860 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_699
timestamp 1649977179
transform 1 0 65412 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_701
timestamp 1649977179
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_713
timestamp 1649977179
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_725
timestamp 1649977179
transform 1 0 67804 0 1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_115_3
timestamp 1649977179
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_15
timestamp 1649977179
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_27
timestamp 1649977179
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_39
timestamp 1649977179
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1649977179
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1649977179
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_115_57
timestamp 1649977179
transform 1 0 6348 0 -1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_115_82
timestamp 1649977179
transform 1 0 8648 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_94
timestamp 1649977179
transform 1 0 9752 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_106
timestamp 1649977179
transform 1 0 10856 0 -1 65280
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_115_113
timestamp 1649977179
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_125
timestamp 1649977179
transform 1 0 12604 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_137
timestamp 1649977179
transform 1 0 13708 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_149
timestamp 1649977179
transform 1 0 14812 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_161
timestamp 1649977179
transform 1 0 15916 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_167
timestamp 1649977179
transform 1 0 16468 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_169
timestamp 1649977179
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_181
timestamp 1649977179
transform 1 0 17756 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_193
timestamp 1649977179
transform 1 0 18860 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_205
timestamp 1649977179
transform 1 0 19964 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_217
timestamp 1649977179
transform 1 0 21068 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_223
timestamp 1649977179
transform 1 0 21620 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_225
timestamp 1649977179
transform 1 0 21804 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_237
timestamp 1649977179
transform 1 0 22908 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_249
timestamp 1649977179
transform 1 0 24012 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_261
timestamp 1649977179
transform 1 0 25116 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_273
timestamp 1649977179
transform 1 0 26220 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_279
timestamp 1649977179
transform 1 0 26772 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_281
timestamp 1649977179
transform 1 0 26956 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_293
timestamp 1649977179
transform 1 0 28060 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_305
timestamp 1649977179
transform 1 0 29164 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_317
timestamp 1649977179
transform 1 0 30268 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_321
timestamp 1649977179
transform 1 0 30636 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_115_325
timestamp 1649977179
transform 1 0 31004 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_332
timestamp 1649977179
transform 1 0 31648 0 -1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_115_358
timestamp 1649977179
transform 1 0 34040 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_370
timestamp 1649977179
transform 1 0 35144 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_382
timestamp 1649977179
transform 1 0 36248 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_115_390
timestamp 1649977179
transform 1 0 36984 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_115_393
timestamp 1649977179
transform 1 0 37260 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_405
timestamp 1649977179
transform 1 0 38364 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_417
timestamp 1649977179
transform 1 0 39468 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_429
timestamp 1649977179
transform 1 0 40572 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_441
timestamp 1649977179
transform 1 0 41676 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_447
timestamp 1649977179
transform 1 0 42228 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_115_449
timestamp 1649977179
transform 1 0 42412 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_115_472
timestamp 1649977179
transform 1 0 44528 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_484
timestamp 1649977179
transform 1 0 45632 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_496
timestamp 1649977179
transform 1 0 46736 0 -1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_115_505
timestamp 1649977179
transform 1 0 47564 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_517
timestamp 1649977179
transform 1 0 48668 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_529
timestamp 1649977179
transform 1 0 49772 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_541
timestamp 1649977179
transform 1 0 50876 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_553
timestamp 1649977179
transform 1 0 51980 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_559
timestamp 1649977179
transform 1 0 52532 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_561
timestamp 1649977179
transform 1 0 52716 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_573
timestamp 1649977179
transform 1 0 53820 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_585
timestamp 1649977179
transform 1 0 54924 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_115_593
timestamp 1649977179
transform 1 0 55660 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_597
timestamp 1649977179
transform 1 0 56028 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_609
timestamp 1649977179
transform 1 0 57132 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_615
timestamp 1649977179
transform 1 0 57684 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_617
timestamp 1649977179
transform 1 0 57868 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_629
timestamp 1649977179
transform 1 0 58972 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_641
timestamp 1649977179
transform 1 0 60076 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_653
timestamp 1649977179
transform 1 0 61180 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_665
timestamp 1649977179
transform 1 0 62284 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_671
timestamp 1649977179
transform 1 0 62836 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_673
timestamp 1649977179
transform 1 0 63020 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_685
timestamp 1649977179
transform 1 0 64124 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_697
timestamp 1649977179
transform 1 0 65228 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_709
timestamp 1649977179
transform 1 0 66332 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_721
timestamp 1649977179
transform 1 0 67436 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_727
timestamp 1649977179
transform 1 0 67988 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_115_729
timestamp 1649977179
transform 1 0 68172 0 -1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1649977179
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1649977179
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1649977179
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1649977179
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_41
timestamp 1649977179
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_53
timestamp 1649977179
transform 1 0 5980 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_116_61
timestamp 1649977179
transform 1 0 6716 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_65
timestamp 1649977179
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_77
timestamp 1649977179
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1649977179
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_85
timestamp 1649977179
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_97
timestamp 1649977179
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_109
timestamp 1649977179
transform 1 0 11132 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_121
timestamp 1649977179
transform 1 0 12236 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_133
timestamp 1649977179
transform 1 0 13340 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_139
timestamp 1649977179
transform 1 0 13892 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_141
timestamp 1649977179
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_153
timestamp 1649977179
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_165
timestamp 1649977179
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_177
timestamp 1649977179
transform 1 0 17388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_189
timestamp 1649977179
transform 1 0 18492 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_195
timestamp 1649977179
transform 1 0 19044 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_197
timestamp 1649977179
transform 1 0 19228 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_209
timestamp 1649977179
transform 1 0 20332 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_221
timestamp 1649977179
transform 1 0 21436 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_233
timestamp 1649977179
transform 1 0 22540 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_245
timestamp 1649977179
transform 1 0 23644 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_251
timestamp 1649977179
transform 1 0 24196 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_253
timestamp 1649977179
transform 1 0 24380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_265
timestamp 1649977179
transform 1 0 25484 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_277
timestamp 1649977179
transform 1 0 26588 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_289
timestamp 1649977179
transform 1 0 27692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_301
timestamp 1649977179
transform 1 0 28796 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_307
timestamp 1649977179
transform 1 0 29348 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_309
timestamp 1649977179
transform 1 0 29532 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_321
timestamp 1649977179
transform 1 0 30636 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_116_329
timestamp 1649977179
transform 1 0 31372 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_116_335
timestamp 1649977179
transform 1 0 31924 0 1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_116_345
timestamp 1649977179
transform 1 0 32844 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_357
timestamp 1649977179
transform 1 0 33948 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_363
timestamp 1649977179
transform 1 0 34500 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_365
timestamp 1649977179
transform 1 0 34684 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_377
timestamp 1649977179
transform 1 0 35788 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_389
timestamp 1649977179
transform 1 0 36892 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_116_400
timestamp 1649977179
transform 1 0 37904 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_412
timestamp 1649977179
transform 1 0 39008 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_116_421
timestamp 1649977179
transform 1 0 39836 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_433
timestamp 1649977179
transform 1 0 40940 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_445
timestamp 1649977179
transform 1 0 42044 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_451
timestamp 1649977179
transform 1 0 42596 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_455
timestamp 1649977179
transform 1 0 42964 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_116_466
timestamp 1649977179
transform 1 0 43976 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_116_474
timestamp 1649977179
transform 1 0 44712 0 1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_116_477
timestamp 1649977179
transform 1 0 44988 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_489
timestamp 1649977179
transform 1 0 46092 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_501
timestamp 1649977179
transform 1 0 47196 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_513
timestamp 1649977179
transform 1 0 48300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_525
timestamp 1649977179
transform 1 0 49404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_531
timestamp 1649977179
transform 1 0 49956 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_533
timestamp 1649977179
transform 1 0 50140 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_545
timestamp 1649977179
transform 1 0 51244 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_557
timestamp 1649977179
transform 1 0 52348 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_569
timestamp 1649977179
transform 1 0 53452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_581
timestamp 1649977179
transform 1 0 54556 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_587
timestamp 1649977179
transform 1 0 55108 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_589
timestamp 1649977179
transform 1 0 55292 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_601
timestamp 1649977179
transform 1 0 56396 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_613
timestamp 1649977179
transform 1 0 57500 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_625
timestamp 1649977179
transform 1 0 58604 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_637
timestamp 1649977179
transform 1 0 59708 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_643
timestamp 1649977179
transform 1 0 60260 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_645
timestamp 1649977179
transform 1 0 60444 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_657
timestamp 1649977179
transform 1 0 61548 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_669
timestamp 1649977179
transform 1 0 62652 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_681
timestamp 1649977179
transform 1 0 63756 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_693
timestamp 1649977179
transform 1 0 64860 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_699
timestamp 1649977179
transform 1 0 65412 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_701
timestamp 1649977179
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_713
timestamp 1649977179
transform 1 0 66700 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_725
timestamp 1649977179
transform 1 0 67804 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1649977179
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1649977179
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_27
timestamp 1649977179
transform 1 0 3588 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_39
timestamp 1649977179
transform 1 0 4692 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_51
timestamp 1649977179
transform 1 0 5796 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_55
timestamp 1649977179
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_57
timestamp 1649977179
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_69
timestamp 1649977179
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_81
timestamp 1649977179
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_93
timestamp 1649977179
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_105
timestamp 1649977179
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_111
timestamp 1649977179
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_113
timestamp 1649977179
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_125
timestamp 1649977179
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_137
timestamp 1649977179
transform 1 0 13708 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_149
timestamp 1649977179
transform 1 0 14812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_161
timestamp 1649977179
transform 1 0 15916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_167
timestamp 1649977179
transform 1 0 16468 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_169
timestamp 1649977179
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_181
timestamp 1649977179
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_193
timestamp 1649977179
transform 1 0 18860 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_205
timestamp 1649977179
transform 1 0 19964 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_217
timestamp 1649977179
transform 1 0 21068 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_223
timestamp 1649977179
transform 1 0 21620 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_225
timestamp 1649977179
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_237
timestamp 1649977179
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_249
timestamp 1649977179
transform 1 0 24012 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_261
timestamp 1649977179
transform 1 0 25116 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_273
timestamp 1649977179
transform 1 0 26220 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_279
timestamp 1649977179
transform 1 0 26772 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_281
timestamp 1649977179
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_293
timestamp 1649977179
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_305
timestamp 1649977179
transform 1 0 29164 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_317
timestamp 1649977179
transform 1 0 30268 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_329
timestamp 1649977179
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_335
timestamp 1649977179
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_337
timestamp 1649977179
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_349
timestamp 1649977179
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_361
timestamp 1649977179
transform 1 0 34316 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_373
timestamp 1649977179
transform 1 0 35420 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_385
timestamp 1649977179
transform 1 0 36524 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_391
timestamp 1649977179
transform 1 0 37076 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_117_393
timestamp 1649977179
transform 1 0 37260 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_416
timestamp 1649977179
transform 1 0 39376 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_428
timestamp 1649977179
transform 1 0 40480 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_440
timestamp 1649977179
transform 1 0 41584 0 -1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_117_449
timestamp 1649977179
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_461
timestamp 1649977179
transform 1 0 43516 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_485
timestamp 1649977179
transform 1 0 45724 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_497
timestamp 1649977179
transform 1 0 46828 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_503
timestamp 1649977179
transform 1 0 47380 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_505
timestamp 1649977179
transform 1 0 47564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_517
timestamp 1649977179
transform 1 0 48668 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_529
timestamp 1649977179
transform 1 0 49772 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_541
timestamp 1649977179
transform 1 0 50876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_553
timestamp 1649977179
transform 1 0 51980 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_559
timestamp 1649977179
transform 1 0 52532 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_561
timestamp 1649977179
transform 1 0 52716 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_573
timestamp 1649977179
transform 1 0 53820 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_585
timestamp 1649977179
transform 1 0 54924 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_597
timestamp 1649977179
transform 1 0 56028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_609
timestamp 1649977179
transform 1 0 57132 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_615
timestamp 1649977179
transform 1 0 57684 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_617
timestamp 1649977179
transform 1 0 57868 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_629
timestamp 1649977179
transform 1 0 58972 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_641
timestamp 1649977179
transform 1 0 60076 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_653
timestamp 1649977179
transform 1 0 61180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_665
timestamp 1649977179
transform 1 0 62284 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_671
timestamp 1649977179
transform 1 0 62836 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_673
timestamp 1649977179
transform 1 0 63020 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_685
timestamp 1649977179
transform 1 0 64124 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_697
timestamp 1649977179
transform 1 0 65228 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_709
timestamp 1649977179
transform 1 0 66332 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_721
timestamp 1649977179
transform 1 0 67436 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_727
timestamp 1649977179
transform 1 0 67988 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_729
timestamp 1649977179
transform 1 0 68172 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1649977179
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1649977179
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1649977179
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1649977179
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_41
timestamp 1649977179
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_53
timestamp 1649977179
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_65
timestamp 1649977179
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1649977179
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1649977179
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_85
timestamp 1649977179
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_97
timestamp 1649977179
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_109
timestamp 1649977179
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_121
timestamp 1649977179
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1649977179
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1649977179
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_141
timestamp 1649977179
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_153
timestamp 1649977179
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_165
timestamp 1649977179
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_177
timestamp 1649977179
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1649977179
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1649977179
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_197
timestamp 1649977179
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_209
timestamp 1649977179
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_221
timestamp 1649977179
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_233
timestamp 1649977179
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_245
timestamp 1649977179
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1649977179
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_253
timestamp 1649977179
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_265
timestamp 1649977179
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_277
timestamp 1649977179
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_289
timestamp 1649977179
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_301
timestamp 1649977179
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_307
timestamp 1649977179
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_309
timestamp 1649977179
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_321
timestamp 1649977179
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_333
timestamp 1649977179
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_345
timestamp 1649977179
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_357
timestamp 1649977179
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_363
timestamp 1649977179
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_365
timestamp 1649977179
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_377
timestamp 1649977179
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_389
timestamp 1649977179
transform 1 0 36892 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_395
timestamp 1649977179
transform 1 0 37444 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_399
timestamp 1649977179
transform 1 0 37812 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_411
timestamp 1649977179
transform 1 0 38916 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1649977179
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_421
timestamp 1649977179
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_433
timestamp 1649977179
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_445
timestamp 1649977179
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_457
timestamp 1649977179
transform 1 0 43148 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_118_468
timestamp 1649977179
transform 1 0 44160 0 1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_118_477
timestamp 1649977179
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_489
timestamp 1649977179
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_501
timestamp 1649977179
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_513
timestamp 1649977179
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_525
timestamp 1649977179
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_531
timestamp 1649977179
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_533
timestamp 1649977179
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_545
timestamp 1649977179
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_557
timestamp 1649977179
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_569
timestamp 1649977179
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_581
timestamp 1649977179
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1649977179
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_589
timestamp 1649977179
transform 1 0 55292 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_601
timestamp 1649977179
transform 1 0 56396 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_613
timestamp 1649977179
transform 1 0 57500 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_625
timestamp 1649977179
transform 1 0 58604 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_637
timestamp 1649977179
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_643
timestamp 1649977179
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_645
timestamp 1649977179
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_657
timestamp 1649977179
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_669
timestamp 1649977179
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_681
timestamp 1649977179
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_693
timestamp 1649977179
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1649977179
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_701
timestamp 1649977179
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_713
timestamp 1649977179
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_725
timestamp 1649977179
transform 1 0 67804 0 1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1649977179
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1649977179
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_27
timestamp 1649977179
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_39
timestamp 1649977179
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1649977179
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1649977179
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_57
timestamp 1649977179
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_69
timestamp 1649977179
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_81
timestamp 1649977179
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_93
timestamp 1649977179
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1649977179
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1649977179
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_113
timestamp 1649977179
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_125
timestamp 1649977179
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_137
timestamp 1649977179
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_149
timestamp 1649977179
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1649977179
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1649977179
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_169
timestamp 1649977179
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_181
timestamp 1649977179
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_193
timestamp 1649977179
transform 1 0 18860 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_205
timestamp 1649977179
transform 1 0 19964 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_217
timestamp 1649977179
transform 1 0 21068 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1649977179
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_225
timestamp 1649977179
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_237
timestamp 1649977179
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_249
timestamp 1649977179
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_261
timestamp 1649977179
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_273
timestamp 1649977179
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1649977179
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_281
timestamp 1649977179
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_293
timestamp 1649977179
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_305
timestamp 1649977179
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_317
timestamp 1649977179
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_329
timestamp 1649977179
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_335
timestamp 1649977179
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_337
timestamp 1649977179
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_349
timestamp 1649977179
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_361
timestamp 1649977179
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_373
timestamp 1649977179
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_385
timestamp 1649977179
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_391
timestamp 1649977179
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_393
timestamp 1649977179
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_405
timestamp 1649977179
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_417
timestamp 1649977179
transform 1 0 39468 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_429
timestamp 1649977179
transform 1 0 40572 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_441
timestamp 1649977179
transform 1 0 41676 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_447
timestamp 1649977179
transform 1 0 42228 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_449
timestamp 1649977179
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_461
timestamp 1649977179
transform 1 0 43516 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_473
timestamp 1649977179
transform 1 0 44620 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_485
timestamp 1649977179
transform 1 0 45724 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_497
timestamp 1649977179
transform 1 0 46828 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1649977179
transform 1 0 47380 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_505
timestamp 1649977179
transform 1 0 47564 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_517
timestamp 1649977179
transform 1 0 48668 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_529
timestamp 1649977179
transform 1 0 49772 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_541
timestamp 1649977179
transform 1 0 50876 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_553
timestamp 1649977179
transform 1 0 51980 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_559
timestamp 1649977179
transform 1 0 52532 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_561
timestamp 1649977179
transform 1 0 52716 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_573
timestamp 1649977179
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_585
timestamp 1649977179
transform 1 0 54924 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_597
timestamp 1649977179
transform 1 0 56028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_609
timestamp 1649977179
transform 1 0 57132 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_615
timestamp 1649977179
transform 1 0 57684 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_617
timestamp 1649977179
transform 1 0 57868 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_629
timestamp 1649977179
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_641
timestamp 1649977179
transform 1 0 60076 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_645
timestamp 1649977179
transform 1 0 60444 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_649
timestamp 1649977179
transform 1 0 60812 0 -1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_119_656
timestamp 1649977179
transform 1 0 61456 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_668
timestamp 1649977179
transform 1 0 62560 0 -1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_119_673
timestamp 1649977179
transform 1 0 63020 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_685
timestamp 1649977179
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_697
timestamp 1649977179
transform 1 0 65228 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_709
timestamp 1649977179
transform 1 0 66332 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_721
timestamp 1649977179
transform 1 0 67436 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_727
timestamp 1649977179
transform 1 0 67988 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_729
timestamp 1649977179
transform 1 0 68172 0 -1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_120_3
timestamp 1649977179
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_15
timestamp 1649977179
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1649977179
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1649977179
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_41
timestamp 1649977179
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_53
timestamp 1649977179
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_65
timestamp 1649977179
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1649977179
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1649977179
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_85
timestamp 1649977179
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_97
timestamp 1649977179
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_109
timestamp 1649977179
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_121
timestamp 1649977179
transform 1 0 12236 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_133
timestamp 1649977179
transform 1 0 13340 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1649977179
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_141
timestamp 1649977179
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_153
timestamp 1649977179
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_165
timestamp 1649977179
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_177
timestamp 1649977179
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_189
timestamp 1649977179
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_195
timestamp 1649977179
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_197
timestamp 1649977179
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_209
timestamp 1649977179
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_221
timestamp 1649977179
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_233
timestamp 1649977179
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1649977179
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1649977179
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_253
timestamp 1649977179
transform 1 0 24380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_265
timestamp 1649977179
transform 1 0 25484 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_277
timestamp 1649977179
transform 1 0 26588 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_289
timestamp 1649977179
transform 1 0 27692 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_301
timestamp 1649977179
transform 1 0 28796 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_307
timestamp 1649977179
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_309
timestamp 1649977179
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_321
timestamp 1649977179
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_333
timestamp 1649977179
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_345
timestamp 1649977179
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_357
timestamp 1649977179
transform 1 0 33948 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1649977179
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_365
timestamp 1649977179
transform 1 0 34684 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_377
timestamp 1649977179
transform 1 0 35788 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_389
timestamp 1649977179
transform 1 0 36892 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_401
timestamp 1649977179
transform 1 0 37996 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_413
timestamp 1649977179
transform 1 0 39100 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_419
timestamp 1649977179
transform 1 0 39652 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_421
timestamp 1649977179
transform 1 0 39836 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_433
timestamp 1649977179
transform 1 0 40940 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_445
timestamp 1649977179
transform 1 0 42044 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_457
timestamp 1649977179
transform 1 0 43148 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_469
timestamp 1649977179
transform 1 0 44252 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_475
timestamp 1649977179
transform 1 0 44804 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_477
timestamp 1649977179
transform 1 0 44988 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_489
timestamp 1649977179
transform 1 0 46092 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_501
timestamp 1649977179
transform 1 0 47196 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_513
timestamp 1649977179
transform 1 0 48300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_525
timestamp 1649977179
transform 1 0 49404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_531
timestamp 1649977179
transform 1 0 49956 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_533
timestamp 1649977179
transform 1 0 50140 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_545
timestamp 1649977179
transform 1 0 51244 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_557
timestamp 1649977179
transform 1 0 52348 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_569
timestamp 1649977179
transform 1 0 53452 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_581
timestamp 1649977179
transform 1 0 54556 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_587
timestamp 1649977179
transform 1 0 55108 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_589
timestamp 1649977179
transform 1 0 55292 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_601
timestamp 1649977179
transform 1 0 56396 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_613
timestamp 1649977179
transform 1 0 57500 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_625
timestamp 1649977179
transform 1 0 58604 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_637
timestamp 1649977179
transform 1 0 59708 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_643
timestamp 1649977179
transform 1 0 60260 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_120_645
timestamp 1649977179
transform 1 0 60444 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_649
timestamp 1649977179
transform 1 0 60812 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_671
timestamp 1649977179
transform 1 0 62836 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_683
timestamp 1649977179
transform 1 0 63940 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_695
timestamp 1649977179
transform 1 0 65044 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_699
timestamp 1649977179
transform 1 0 65412 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_701
timestamp 1649977179
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_713
timestamp 1649977179
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_725
timestamp 1649977179
transform 1 0 67804 0 1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1649977179
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1649977179
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_27
timestamp 1649977179
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_39
timestamp 1649977179
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1649977179
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1649977179
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_57
timestamp 1649977179
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_69
timestamp 1649977179
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_81
timestamp 1649977179
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_93
timestamp 1649977179
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1649977179
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1649977179
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_113
timestamp 1649977179
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_125
timestamp 1649977179
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_137
timestamp 1649977179
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_149
timestamp 1649977179
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1649977179
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1649977179
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_169
timestamp 1649977179
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_181
timestamp 1649977179
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_193
timestamp 1649977179
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_205
timestamp 1649977179
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_217
timestamp 1649977179
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_223
timestamp 1649977179
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_225
timestamp 1649977179
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_237
timestamp 1649977179
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_249
timestamp 1649977179
transform 1 0 24012 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_261
timestamp 1649977179
transform 1 0 25116 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_273
timestamp 1649977179
transform 1 0 26220 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1649977179
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_281
timestamp 1649977179
transform 1 0 26956 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_293
timestamp 1649977179
transform 1 0 28060 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_305
timestamp 1649977179
transform 1 0 29164 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_317
timestamp 1649977179
transform 1 0 30268 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_329
timestamp 1649977179
transform 1 0 31372 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_335
timestamp 1649977179
transform 1 0 31924 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_337
timestamp 1649977179
transform 1 0 32108 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_349
timestamp 1649977179
transform 1 0 33212 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_361
timestamp 1649977179
transform 1 0 34316 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_373
timestamp 1649977179
transform 1 0 35420 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_385
timestamp 1649977179
transform 1 0 36524 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_391
timestamp 1649977179
transform 1 0 37076 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_393
timestamp 1649977179
transform 1 0 37260 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_405
timestamp 1649977179
transform 1 0 38364 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_417
timestamp 1649977179
transform 1 0 39468 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_429
timestamp 1649977179
transform 1 0 40572 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_441
timestamp 1649977179
transform 1 0 41676 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_447
timestamp 1649977179
transform 1 0 42228 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_449
timestamp 1649977179
transform 1 0 42412 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_461
timestamp 1649977179
transform 1 0 43516 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_473
timestamp 1649977179
transform 1 0 44620 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_485
timestamp 1649977179
transform 1 0 45724 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_497
timestamp 1649977179
transform 1 0 46828 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_503
timestamp 1649977179
transform 1 0 47380 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_505
timestamp 1649977179
transform 1 0 47564 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_517
timestamp 1649977179
transform 1 0 48668 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_529
timestamp 1649977179
transform 1 0 49772 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_541
timestamp 1649977179
transform 1 0 50876 0 -1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_121_546
timestamp 1649977179
transform 1 0 51336 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_558
timestamp 1649977179
transform 1 0 52440 0 -1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_121_561
timestamp 1649977179
transform 1 0 52716 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_573
timestamp 1649977179
transform 1 0 53820 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_585
timestamp 1649977179
transform 1 0 54924 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_121_597
timestamp 1649977179
transform 1 0 56028 0 -1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_121_603
timestamp 1649977179
transform 1 0 56580 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_121_615
timestamp 1649977179
transform 1 0 57684 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_617
timestamp 1649977179
transform 1 0 57868 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_650
timestamp 1649977179
transform 1 0 60904 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_662
timestamp 1649977179
transform 1 0 62008 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_121_670
timestamp 1649977179
transform 1 0 62744 0 -1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_121_673
timestamp 1649977179
transform 1 0 63020 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_685
timestamp 1649977179
transform 1 0 64124 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_697
timestamp 1649977179
transform 1 0 65228 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_709
timestamp 1649977179
transform 1 0 66332 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_721
timestamp 1649977179
transform 1 0 67436 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_727
timestamp 1649977179
transform 1 0 67988 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_121_729
timestamp 1649977179
transform 1 0 68172 0 -1 68544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_122_3
timestamp 1649977179
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_15
timestamp 1649977179
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1649977179
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1649977179
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_41
timestamp 1649977179
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_53
timestamp 1649977179
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_65
timestamp 1649977179
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1649977179
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1649977179
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_85
timestamp 1649977179
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_97
timestamp 1649977179
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_109
timestamp 1649977179
transform 1 0 11132 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_121
timestamp 1649977179
transform 1 0 12236 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_133
timestamp 1649977179
transform 1 0 13340 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_139
timestamp 1649977179
transform 1 0 13892 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_141
timestamp 1649977179
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_153
timestamp 1649977179
transform 1 0 15180 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_165
timestamp 1649977179
transform 1 0 16284 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_177
timestamp 1649977179
transform 1 0 17388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_189
timestamp 1649977179
transform 1 0 18492 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_195
timestamp 1649977179
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_197
timestamp 1649977179
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_209
timestamp 1649977179
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_221
timestamp 1649977179
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_233
timestamp 1649977179
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_245
timestamp 1649977179
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_251
timestamp 1649977179
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_253
timestamp 1649977179
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_265
timestamp 1649977179
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_277
timestamp 1649977179
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_289
timestamp 1649977179
transform 1 0 27692 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_301
timestamp 1649977179
transform 1 0 28796 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_307
timestamp 1649977179
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_309
timestamp 1649977179
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_321
timestamp 1649977179
transform 1 0 30636 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_333
timestamp 1649977179
transform 1 0 31740 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_345
timestamp 1649977179
transform 1 0 32844 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_357
timestamp 1649977179
transform 1 0 33948 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_363
timestamp 1649977179
transform 1 0 34500 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_365
timestamp 1649977179
transform 1 0 34684 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_377
timestamp 1649977179
transform 1 0 35788 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_389
timestamp 1649977179
transform 1 0 36892 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_401
timestamp 1649977179
transform 1 0 37996 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_413
timestamp 1649977179
transform 1 0 39100 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_419
timestamp 1649977179
transform 1 0 39652 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_421
timestamp 1649977179
transform 1 0 39836 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_433
timestamp 1649977179
transform 1 0 40940 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_445
timestamp 1649977179
transform 1 0 42044 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_457
timestamp 1649977179
transform 1 0 43148 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_469
timestamp 1649977179
transform 1 0 44252 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_475
timestamp 1649977179
transform 1 0 44804 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_477
timestamp 1649977179
transform 1 0 44988 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_489
timestamp 1649977179
transform 1 0 46092 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_514
timestamp 1649977179
transform 1 0 48392 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_122_521
timestamp 1649977179
transform 1 0 49036 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_529
timestamp 1649977179
transform 1 0 49772 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_122_533
timestamp 1649977179
transform 1 0 50140 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_541
timestamp 1649977179
transform 1 0 50876 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_563
timestamp 1649977179
transform 1 0 52900 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_575
timestamp 1649977179
transform 1 0 54004 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_587
timestamp 1649977179
transform 1 0 55108 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_589
timestamp 1649977179
transform 1 0 55292 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_122_597
timestamp 1649977179
transform 1 0 56028 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_122_620
timestamp 1649977179
transform 1 0 58144 0 1 68544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_122_631
timestamp 1649977179
transform 1 0 59156 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_643
timestamp 1649977179
transform 1 0 60260 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_645
timestamp 1649977179
transform 1 0 60444 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_657
timestamp 1649977179
transform 1 0 61548 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_669
timestamp 1649977179
transform 1 0 62652 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_681
timestamp 1649977179
transform 1 0 63756 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_693
timestamp 1649977179
transform 1 0 64860 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_699
timestamp 1649977179
transform 1 0 65412 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_701
timestamp 1649977179
transform 1 0 65596 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_713
timestamp 1649977179
transform 1 0 66700 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_725
timestamp 1649977179
transform 1 0 67804 0 1 68544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_123_12
timestamp 1649977179
transform 1 0 2208 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_24
timestamp 1649977179
transform 1 0 3312 0 -1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_123_29
timestamp 1649977179
transform 1 0 3772 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_41
timestamp 1649977179
transform 1 0 4876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_53
timestamp 1649977179
transform 1 0 5980 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_57
timestamp 1649977179
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_69
timestamp 1649977179
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_81
timestamp 1649977179
transform 1 0 8556 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_85
timestamp 1649977179
transform 1 0 8924 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_97
timestamp 1649977179
transform 1 0 10028 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_109
timestamp 1649977179
transform 1 0 11132 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_113
timestamp 1649977179
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_125
timestamp 1649977179
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_137
timestamp 1649977179
transform 1 0 13708 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_141
timestamp 1649977179
transform 1 0 14076 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_153
timestamp 1649977179
transform 1 0 15180 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_165
timestamp 1649977179
transform 1 0 16284 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_169
timestamp 1649977179
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_181
timestamp 1649977179
transform 1 0 17756 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_193
timestamp 1649977179
transform 1 0 18860 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_197
timestamp 1649977179
transform 1 0 19228 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_209
timestamp 1649977179
transform 1 0 20332 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_221
timestamp 1649977179
transform 1 0 21436 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_225
timestamp 1649977179
transform 1 0 21804 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_237
timestamp 1649977179
transform 1 0 22908 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_249
timestamp 1649977179
transform 1 0 24012 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_253
timestamp 1649977179
transform 1 0 24380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_265
timestamp 1649977179
transform 1 0 25484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_277
timestamp 1649977179
transform 1 0 26588 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_281
timestamp 1649977179
transform 1 0 26956 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_293
timestamp 1649977179
transform 1 0 28060 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_305
timestamp 1649977179
transform 1 0 29164 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_309
timestamp 1649977179
transform 1 0 29532 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_321
timestamp 1649977179
transform 1 0 30636 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_333
timestamp 1649977179
transform 1 0 31740 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_337
timestamp 1649977179
transform 1 0 32108 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_349
timestamp 1649977179
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_361
timestamp 1649977179
transform 1 0 34316 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_365
timestamp 1649977179
transform 1 0 34684 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_377
timestamp 1649977179
transform 1 0 35788 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_389
timestamp 1649977179
transform 1 0 36892 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_393
timestamp 1649977179
transform 1 0 37260 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_405
timestamp 1649977179
transform 1 0 38364 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_417
timestamp 1649977179
transform 1 0 39468 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_421
timestamp 1649977179
transform 1 0 39836 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_433
timestamp 1649977179
transform 1 0 40940 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_445
timestamp 1649977179
transform 1 0 42044 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_449
timestamp 1649977179
transform 1 0 42412 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_461
timestamp 1649977179
transform 1 0 43516 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_473
timestamp 1649977179
transform 1 0 44620 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_477
timestamp 1649977179
transform 1 0 44988 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_489
timestamp 1649977179
transform 1 0 46092 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_493
timestamp 1649977179
transform 1 0 46460 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_123_497
timestamp 1649977179
transform 1 0 46828 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_503
timestamp 1649977179
transform 1 0 47380 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_505
timestamp 1649977179
transform 1 0 47564 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_517
timestamp 1649977179
transform 1 0 48668 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_529
timestamp 1649977179
transform 1 0 49772 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_123_533
timestamp 1649977179
transform 1 0 50140 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_123_541
timestamp 1649977179
transform 1 0 50876 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_123_546
timestamp 1649977179
transform 1 0 51336 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_558
timestamp 1649977179
transform 1 0 52440 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_123_561
timestamp 1649977179
transform 1 0 52716 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_573
timestamp 1649977179
transform 1 0 53820 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_585
timestamp 1649977179
transform 1 0 54924 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_123_589
timestamp 1649977179
transform 1 0 55292 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_123_601
timestamp 1649977179
transform 1 0 56396 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_123_608
timestamp 1649977179
transform 1 0 57040 0 -1 69632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_123_617
timestamp 1649977179
transform 1 0 57868 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_123_629
timestamp 1649977179
transform 1 0 58972 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_633
timestamp 1649977179
transform 1 0 59340 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_123_641
timestamp 1649977179
transform 1 0 60076 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_645
timestamp 1649977179
transform 1 0 60444 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_657
timestamp 1649977179
transform 1 0 61548 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_669
timestamp 1649977179
transform 1 0 62652 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_673
timestamp 1649977179
transform 1 0 63020 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_685
timestamp 1649977179
transform 1 0 64124 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_697
timestamp 1649977179
transform 1 0 65228 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_701
timestamp 1649977179
transform 1 0 65596 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_713
timestamp 1649977179
transform 1 0 66700 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_719
timestamp 1649977179
transform 1 0 67252 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_123_724
timestamp 1649977179
transform 1 0 67712 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_729
timestamp 1649977179
transform 1 0 68172 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 68816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 68816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 68816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 68816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 68816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 68816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 68816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 68816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 68816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 68816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 68816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 68816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 68816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 68816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 68816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 68816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 68816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 68816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 68816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 68816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 68816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 68816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 68816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 68816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 68816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 68816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 68816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 68816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 68816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 68816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 68816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 68816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 68816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 68816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 68816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 68816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 68816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 68816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 68816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 68816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 68816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 68816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 68816 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 68816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 68816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 68816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 68816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 68816 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 68816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 68816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 68816 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 68816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 68816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 68816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 68816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 68816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 68816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 68816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 68816 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 68816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 68816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 68816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 68816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 68816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 68816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 68816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 68816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 68816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 68816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 68816 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 68816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 68816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 68816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 68816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 68816 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 68816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 68816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 68816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 68816 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 68816 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 68816 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 68816 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 68816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 68816 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 68816 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 68816 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 68816 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 68816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 68816 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 68816 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 68816 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 68816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 68816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 68816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 68816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1649977179
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1649977179
transform -1 0 68816 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1649977179
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1649977179
transform -1 0 68816 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1649977179
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1649977179
transform -1 0 68816 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1649977179
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1649977179
transform -1 0 68816 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1649977179
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1649977179
transform -1 0 68816 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1649977179
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1649977179
transform -1 0 68816 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1649977179
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1649977179
transform -1 0 68816 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1649977179
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1649977179
transform -1 0 68816 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1649977179
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1649977179
transform -1 0 68816 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1649977179
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1649977179
transform -1 0 68816 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1649977179
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1649977179
transform -1 0 68816 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1649977179
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1649977179
transform -1 0 68816 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1649977179
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1649977179
transform -1 0 68816 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1649977179
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1649977179
transform -1 0 68816 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1649977179
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1649977179
transform -1 0 68816 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1649977179
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1649977179
transform -1 0 68816 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1649977179
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1649977179
transform -1 0 68816 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1649977179
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1649977179
transform -1 0 68816 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1649977179
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1649977179
transform -1 0 68816 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1649977179
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1649977179
transform -1 0 68816 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1649977179
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1649977179
transform -1 0 68816 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1649977179
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1649977179
transform -1 0 68816 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1649977179
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1649977179
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1649977179
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1649977179
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1649977179
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1649977179
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1649977179
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1649977179
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1649977179
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1649977179
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1649977179
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1649977179
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1649977179
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1649977179
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1649977179
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1649977179
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1649977179
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1649977179
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1649977179
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1649977179
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1649977179
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1649977179
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1649977179
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1649977179
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1649977179
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1649977179
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1649977179
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1649977179
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1649977179
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1649977179
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1649977179
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1649977179
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1649977179
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1649977179
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1649977179
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1649977179
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1649977179
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1649977179
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1649977179
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1649977179
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1649977179
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1649977179
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1649977179
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1649977179
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1649977179
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1649977179
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1649977179
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1649977179
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1649977179
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1649977179
transform 1 0 60352 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1649977179
transform 1 0 65504 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1649977179
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1649977179
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1649977179
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1649977179
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1649977179
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1649977179
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1649977179
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1649977179
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1649977179
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1649977179
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1649977179
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1649977179
transform 1 0 62928 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1649977179
transform 1 0 68080 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1649977179
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1649977179
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1649977179
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1649977179
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1649977179
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1649977179
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1649977179
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1649977179
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1649977179
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1649977179
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1649977179
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1649977179
transform 1 0 60352 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1649977179
transform 1 0 65504 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1649977179
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1649977179
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1649977179
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1649977179
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1649977179
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1649977179
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1649977179
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1649977179
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1649977179
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1649977179
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1649977179
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1649977179
transform 1 0 62928 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1649977179
transform 1 0 68080 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1649977179
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1649977179
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1649977179
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1649977179
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1649977179
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1649977179
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1649977179
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1649977179
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1649977179
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1649977179
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1649977179
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1649977179
transform 1 0 60352 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1649977179
transform 1 0 65504 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1649977179
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1649977179
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1649977179
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1649977179
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1649977179
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1649977179
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1649977179
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1649977179
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1660
timestamp 1649977179
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1661
timestamp 1649977179
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1662
timestamp 1649977179
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1663
timestamp 1649977179
transform 1 0 62928 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1664
timestamp 1649977179
transform 1 0 68080 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1665
timestamp 1649977179
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1666
timestamp 1649977179
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1667
timestamp 1649977179
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1668
timestamp 1649977179
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1669
timestamp 1649977179
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1670
timestamp 1649977179
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1671
timestamp 1649977179
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1672
timestamp 1649977179
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1673
timestamp 1649977179
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1674
timestamp 1649977179
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1675
timestamp 1649977179
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1676
timestamp 1649977179
transform 1 0 60352 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1677
timestamp 1649977179
transform 1 0 65504 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1678
timestamp 1649977179
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1679
timestamp 1649977179
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1680
timestamp 1649977179
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1681
timestamp 1649977179
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1682
timestamp 1649977179
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1683
timestamp 1649977179
transform 1 0 32016 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1684
timestamp 1649977179
transform 1 0 37168 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1685
timestamp 1649977179
transform 1 0 42320 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1686
timestamp 1649977179
transform 1 0 47472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1687
timestamp 1649977179
transform 1 0 52624 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1688
timestamp 1649977179
transform 1 0 57776 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1689
timestamp 1649977179
transform 1 0 62928 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1690
timestamp 1649977179
transform 1 0 68080 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1691
timestamp 1649977179
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1692
timestamp 1649977179
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1693
timestamp 1649977179
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1694
timestamp 1649977179
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1695
timestamp 1649977179
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1696
timestamp 1649977179
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1697
timestamp 1649977179
transform 1 0 34592 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1698
timestamp 1649977179
transform 1 0 39744 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1699
timestamp 1649977179
transform 1 0 44896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1700
timestamp 1649977179
transform 1 0 50048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1701
timestamp 1649977179
transform 1 0 55200 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1702
timestamp 1649977179
transform 1 0 60352 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1703
timestamp 1649977179
transform 1 0 65504 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1704
timestamp 1649977179
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1705
timestamp 1649977179
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1706
timestamp 1649977179
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1707
timestamp 1649977179
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1708
timestamp 1649977179
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1709
timestamp 1649977179
transform 1 0 32016 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1710
timestamp 1649977179
transform 1 0 37168 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1711
timestamp 1649977179
transform 1 0 42320 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1712
timestamp 1649977179
transform 1 0 47472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1713
timestamp 1649977179
transform 1 0 52624 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1714
timestamp 1649977179
transform 1 0 57776 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1715
timestamp 1649977179
transform 1 0 62928 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1716
timestamp 1649977179
transform 1 0 68080 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1717
timestamp 1649977179
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1718
timestamp 1649977179
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1719
timestamp 1649977179
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1720
timestamp 1649977179
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1721
timestamp 1649977179
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1722
timestamp 1649977179
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1723
timestamp 1649977179
transform 1 0 34592 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1724
timestamp 1649977179
transform 1 0 39744 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1725
timestamp 1649977179
transform 1 0 44896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1726
timestamp 1649977179
transform 1 0 50048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1727
timestamp 1649977179
transform 1 0 55200 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1728
timestamp 1649977179
transform 1 0 60352 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1729
timestamp 1649977179
transform 1 0 65504 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1730
timestamp 1649977179
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1731
timestamp 1649977179
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1732
timestamp 1649977179
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1733
timestamp 1649977179
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1734
timestamp 1649977179
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1735
timestamp 1649977179
transform 1 0 32016 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1736
timestamp 1649977179
transform 1 0 37168 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1737
timestamp 1649977179
transform 1 0 42320 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1738
timestamp 1649977179
transform 1 0 47472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1739
timestamp 1649977179
transform 1 0 52624 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1740
timestamp 1649977179
transform 1 0 57776 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1741
timestamp 1649977179
transform 1 0 62928 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1742
timestamp 1649977179
transform 1 0 68080 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1743
timestamp 1649977179
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1744
timestamp 1649977179
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1745
timestamp 1649977179
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1746
timestamp 1649977179
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1747
timestamp 1649977179
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1748
timestamp 1649977179
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1749
timestamp 1649977179
transform 1 0 34592 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1750
timestamp 1649977179
transform 1 0 39744 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1751
timestamp 1649977179
transform 1 0 44896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1752
timestamp 1649977179
transform 1 0 50048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1753
timestamp 1649977179
transform 1 0 55200 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1754
timestamp 1649977179
transform 1 0 60352 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1755
timestamp 1649977179
transform 1 0 65504 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1756
timestamp 1649977179
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1757
timestamp 1649977179
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1758
timestamp 1649977179
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1759
timestamp 1649977179
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1760
timestamp 1649977179
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1761
timestamp 1649977179
transform 1 0 32016 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1762
timestamp 1649977179
transform 1 0 37168 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1763
timestamp 1649977179
transform 1 0 42320 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1764
timestamp 1649977179
transform 1 0 47472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1765
timestamp 1649977179
transform 1 0 52624 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1766
timestamp 1649977179
transform 1 0 57776 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1767
timestamp 1649977179
transform 1 0 62928 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1768
timestamp 1649977179
transform 1 0 68080 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1769
timestamp 1649977179
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1770
timestamp 1649977179
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1771
timestamp 1649977179
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1772
timestamp 1649977179
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1773
timestamp 1649977179
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1774
timestamp 1649977179
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1775
timestamp 1649977179
transform 1 0 34592 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1776
timestamp 1649977179
transform 1 0 39744 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1777
timestamp 1649977179
transform 1 0 44896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1778
timestamp 1649977179
transform 1 0 50048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1779
timestamp 1649977179
transform 1 0 55200 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1780
timestamp 1649977179
transform 1 0 60352 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1781
timestamp 1649977179
transform 1 0 65504 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1782
timestamp 1649977179
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1783
timestamp 1649977179
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1784
timestamp 1649977179
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1785
timestamp 1649977179
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1786
timestamp 1649977179
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1787
timestamp 1649977179
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1788
timestamp 1649977179
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1789
timestamp 1649977179
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1790
timestamp 1649977179
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1791
timestamp 1649977179
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1792
timestamp 1649977179
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1793
timestamp 1649977179
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1794
timestamp 1649977179
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1795
timestamp 1649977179
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1796
timestamp 1649977179
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1797
timestamp 1649977179
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1798
timestamp 1649977179
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1799
timestamp 1649977179
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1800
timestamp 1649977179
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1801
timestamp 1649977179
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1802
timestamp 1649977179
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1803
timestamp 1649977179
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1804
timestamp 1649977179
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1805
timestamp 1649977179
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1806
timestamp 1649977179
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1807
timestamp 1649977179
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1808
timestamp 1649977179
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1809
timestamp 1649977179
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1810
timestamp 1649977179
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1811
timestamp 1649977179
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1812
timestamp 1649977179
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1813
timestamp 1649977179
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1814
timestamp 1649977179
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1815
timestamp 1649977179
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1816
timestamp 1649977179
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1817
timestamp 1649977179
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1818
timestamp 1649977179
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1819
timestamp 1649977179
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1820
timestamp 1649977179
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1821
timestamp 1649977179
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1822
timestamp 1649977179
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1823
timestamp 1649977179
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1824
timestamp 1649977179
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1825
timestamp 1649977179
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1826
timestamp 1649977179
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1827
timestamp 1649977179
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1828
timestamp 1649977179
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1829
timestamp 1649977179
transform 1 0 44896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1830
timestamp 1649977179
transform 1 0 50048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1831
timestamp 1649977179
transform 1 0 55200 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1832
timestamp 1649977179
transform 1 0 60352 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1833
timestamp 1649977179
transform 1 0 65504 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1834
timestamp 1649977179
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1835
timestamp 1649977179
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1836
timestamp 1649977179
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1837
timestamp 1649977179
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1838
timestamp 1649977179
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1839
timestamp 1649977179
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1840
timestamp 1649977179
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1841
timestamp 1649977179
transform 1 0 42320 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1842
timestamp 1649977179
transform 1 0 47472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1843
timestamp 1649977179
transform 1 0 52624 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1844
timestamp 1649977179
transform 1 0 57776 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1845
timestamp 1649977179
transform 1 0 62928 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1846
timestamp 1649977179
transform 1 0 68080 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1847
timestamp 1649977179
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1848
timestamp 1649977179
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1849
timestamp 1649977179
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1850
timestamp 1649977179
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1851
timestamp 1649977179
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1852
timestamp 1649977179
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1853
timestamp 1649977179
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1854
timestamp 1649977179
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1855
timestamp 1649977179
transform 1 0 44896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1856
timestamp 1649977179
transform 1 0 50048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1857
timestamp 1649977179
transform 1 0 55200 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1858
timestamp 1649977179
transform 1 0 60352 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1859
timestamp 1649977179
transform 1 0 65504 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1860
timestamp 1649977179
transform 1 0 3680 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1861
timestamp 1649977179
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1862
timestamp 1649977179
transform 1 0 8832 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1863
timestamp 1649977179
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1864
timestamp 1649977179
transform 1 0 13984 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1865
timestamp 1649977179
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1866
timestamp 1649977179
transform 1 0 19136 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1867
timestamp 1649977179
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1868
timestamp 1649977179
transform 1 0 24288 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1869
timestamp 1649977179
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1870
timestamp 1649977179
transform 1 0 29440 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1871
timestamp 1649977179
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1872
timestamp 1649977179
transform 1 0 34592 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1873
timestamp 1649977179
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1874
timestamp 1649977179
transform 1 0 39744 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1875
timestamp 1649977179
transform 1 0 42320 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1876
timestamp 1649977179
transform 1 0 44896 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1877
timestamp 1649977179
transform 1 0 47472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1878
timestamp 1649977179
transform 1 0 50048 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1879
timestamp 1649977179
transform 1 0 52624 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1880
timestamp 1649977179
transform 1 0 55200 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1881
timestamp 1649977179
transform 1 0 57776 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1882
timestamp 1649977179
transform 1 0 60352 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1883
timestamp 1649977179
transform 1 0 62928 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1884
timestamp 1649977179
transform 1 0 65504 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1885
timestamp 1649977179
transform 1 0 68080 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _244_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31372 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _245_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43976 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _246_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 44068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _247_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1649977179
transform 1 0 26128 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1649977179
transform 1 0 26404 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1649977179
transform 1 0 9476 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1649977179
transform 1 0 8096 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _253_
timestamp 1649977179
transform 1 0 37720 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1649977179
transform 1 0 27048 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1649977179
transform 1 0 23460 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1649977179
transform 1 0 50140 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1649977179
transform 1 0 54464 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1649977179
transform 1 0 52072 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _259_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43608 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  _260_
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1649977179
transform 1 0 53176 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1649977179
transform 1 0 51244 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1649977179
transform 1 0 26864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1649977179
transform 1 0 25024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _266_
timestamp 1649977179
transform 1 0 44160 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1649977179
transform 1 0 32292 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1649977179
transform 1 0 33120 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1649977179
transform 1 0 54372 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _272_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 45080 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1649977179
transform 1 0 64492 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1649977179
transform 1 0 57868 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1649977179
transform 1 0 64676 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1649977179
transform 1 0 64952 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _278_
timestamp 1649977179
transform 1 0 43700 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1649977179
transform 1 0 43700 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1649977179
transform 1 0 42688 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1649977179
transform 1 0 37352 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1649977179
transform 1 0 37628 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1649977179
transform 1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _284_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1649977179
transform 1 0 32384 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1649977179
transform 1 0 62652 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1649977179
transform 1 0 63112 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1649977179
transform 1 0 27784 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1649977179
transform 1 0 62928 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _290_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20516 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _291_
timestamp 1649977179
transform 1 0 20608 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1649977179
transform 1 0 34776 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1649977179
transform 1 0 9752 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1649977179
transform 1 0 10764 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1649977179
transform 1 0 34684 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _297_
timestamp 1649977179
transform 1 0 20608 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1649977179
transform 1 0 38180 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1649977179
transform 1 0 4968 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1649977179
transform 1 0 35236 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1649977179
transform 1 0 5428 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1649977179
transform 1 0 5612 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _303_
timestamp 1649977179
transform 1 0 21528 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1649977179
transform 1 0 36800 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1649977179
transform 1 0 19872 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1649977179
transform 1 0 35512 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1649977179
transform 1 0 28520 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1649977179
transform 1 0 22080 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _309_
timestamp 1649977179
transform 1 0 19688 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1649977179
transform 1 0 21344 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1649977179
transform 1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1649977179
transform 1 0 4968 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1649977179
transform 1 0 12788 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1649977179
transform 1 0 5428 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _315_
timestamp 1649977179
transform 1 0 20516 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1649977179
transform 1 0 30636 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1649977179
transform 1 0 28612 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1649977179
transform 1 0 6992 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1649977179
transform 1 0 6624 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1649977179
transform 1 0 7176 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _321_
timestamp 1649977179
transform 1 0 42136 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  _322_
timestamp 1649977179
transform 1 0 42320 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1649977179
transform 1 0 43332 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1649977179
transform 1 0 22540 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1649977179
transform 1 0 54372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1649977179
transform 1 0 51152 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _328_
timestamp 1649977179
transform 1 0 42412 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1649977179
transform 1 0 56948 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1649977179
transform 1 0 42320 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1649977179
transform 1 0 58972 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1649977179
transform 1 0 47564 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1649977179
transform 1 0 48484 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _334_
timestamp 1649977179
transform 1 0 42780 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1649977179
transform 1 0 41676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1649977179
transform 1 0 43424 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1649977179
transform 1 0 27048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _340_
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1649977179
transform 1 0 57868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1649977179
transform 1 0 50508 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1649977179
transform 1 0 46552 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1649977179
transform 1 0 55568 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _346_
timestamp 1649977179
transform 1 0 41400 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1649977179
transform 1 0 44068 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1649977179
transform 1 0 51060 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1649977179
transform 1 0 54188 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1649977179
transform 1 0 30268 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _352_
timestamp 1649977179
transform 1 0 47656 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1649977179
transform 1 0 28796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1649977179
transform 1 0 60720 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1649977179
transform 1 0 61824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1649977179
transform 1 0 33396 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1649977179
transform 1 0 60352 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _358_
timestamp 1649977179
transform 1 0 48760 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1649977179
transform 1 0 30544 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1649977179
transform 1 0 63204 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1649977179
transform 1 0 63664 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1649977179
transform 1 0 63388 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1649977179
transform 1 0 35144 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _364_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 48944 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1649977179
transform 1 0 58880 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1649977179
transform 1 0 51060 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1649977179
transform 1 0 60536 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1649977179
transform 1 0 56304 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1649977179
transform 1 0 48760 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _370_
timestamp 1649977179
transform 1 0 49404 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1649977179
transform 1 0 67436 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1649977179
transform 1 0 67068 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1649977179
transform 1 0 67436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1649977179
transform 1 0 45908 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1649977179
transform 1 0 67436 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1649977179
transform 1 0 43516 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1649977179
transform 1 0 14996 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1649977179
transform 1 0 12604 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _379_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33948 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _380_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 31280 0 1 64192
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _381_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31280 0 1 63104
box -38 -48 1510 592
use sky130_fd_sc_hd__ebufn_8  _489_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32568 0 -1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _490__6 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _490_
timestamp 1649977179
transform 1 0 12144 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _491__7
timestamp 1649977179
transform 1 0 51152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _491_
timestamp 1649977179
transform 1 0 50324 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _492__8
timestamp 1649977179
transform 1 0 58236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _492_
timestamp 1649977179
transform 1 0 58144 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _493__9
timestamp 1649977179
transform 1 0 27692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _493_
timestamp 1649977179
transform 1 0 27600 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _494_
timestamp 1649977179
transform 1 0 26864 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _494__10
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _495_
timestamp 1649977179
transform 1 0 39376 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _495__11
timestamp 1649977179
transform 1 0 38732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _496__12
timestamp 1649977179
transform 1 0 43332 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _496_
timestamp 1649977179
transform 1 0 42872 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _497_
timestamp 1649977179
transform 1 0 40664 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _497__13
timestamp 1649977179
transform 1 0 40664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _498__14
timestamp 1649977179
transform 1 0 48484 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _498_
timestamp 1649977179
transform 1 0 48392 0 -1 57664
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _499__15
timestamp 1649977179
transform 1 0 46460 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _499_
timestamp 1649977179
transform 1 0 47104 0 1 59840
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _500__16
timestamp 1649977179
transform 1 0 59616 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _500_
timestamp 1649977179
transform 1 0 59616 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _501__17
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _501_
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _502__18
timestamp 1649977179
transform 1 0 57132 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _502_
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _503__19
timestamp 1649977179
transform 1 0 51336 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _503_
timestamp 1649977179
transform 1 0 51336 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _504__20
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _504_
timestamp 1649977179
transform 1 0 54740 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _505__21
timestamp 1649977179
transform 1 0 60536 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _505_
timestamp 1649977179
transform 1 0 60444 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _506_
timestamp 1649977179
transform 1 0 32292 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _506__22
timestamp 1649977179
transform 1 0 32752 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _507__23
timestamp 1649977179
transform 1 0 22908 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _507_
timestamp 1649977179
transform 1 0 21988 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _508_
timestamp 1649977179
transform 1 0 43240 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _508__24
timestamp 1649977179
transform 1 0 43332 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _509__25
timestamp 1649977179
transform 1 0 25760 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _509_
timestamp 1649977179
transform 1 0 26404 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _510__26
timestamp 1649977179
transform 1 0 6992 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _510_
timestamp 1649977179
transform 1 0 6900 0 -1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _511__27
timestamp 1649977179
transform 1 0 6808 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _511_
timestamp 1649977179
transform 1 0 6716 0 -1 65280
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _512__28
timestamp 1649977179
transform 1 0 29532 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _512_
timestamp 1649977179
transform 1 0 29256 0 -1 64192
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _513__29
timestamp 1649977179
transform 1 0 5244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _513_
timestamp 1649977179
transform 1 0 5244 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _514__30
timestamp 1649977179
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _514_
timestamp 1649977179
transform 1 0 12788 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _515__31
timestamp 1649977179
transform 1 0 5244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _515_
timestamp 1649977179
transform 1 0 5152 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _516__32
timestamp 1649977179
transform 1 0 22264 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _516_
timestamp 1649977179
transform 1 0 22264 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _517__33
timestamp 1649977179
transform 1 0 28520 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _517_
timestamp 1649977179
transform 1 0 27416 0 -1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _518__34
timestamp 1649977179
transform 1 0 35512 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _518_
timestamp 1649977179
transform 1 0 35420 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _519__35
timestamp 1649977179
transform 1 0 37168 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _519_
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _520__36
timestamp 1649977179
transform 1 0 5336 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _520_
timestamp 1649977179
transform 1 0 5244 0 1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _521__37
timestamp 1649977179
transform 1 0 35328 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _521_
timestamp 1649977179
transform 1 0 34868 0 -1 51136
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _522__38
timestamp 1649977179
transform 1 0 14720 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _522_
timestamp 1649977179
transform 1 0 14720 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _523_
timestamp 1649977179
transform 1 0 5612 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _523__39
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _524_
timestamp 1649977179
transform 1 0 34868 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _524__40
timestamp 1649977179
transform 1 0 34960 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _525__41
timestamp 1649977179
transform 1 0 11408 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _525_
timestamp 1649977179
transform 1 0 10580 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _526__42
timestamp 1649977179
transform 1 0 9568 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _526_
timestamp 1649977179
transform 1 0 9568 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _527__43
timestamp 1649977179
transform 1 0 35144 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _527_
timestamp 1649977179
transform 1 0 35052 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _528__44
timestamp 1649977179
transform 1 0 62192 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _528_
timestamp 1649977179
transform 1 0 62192 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _529__45
timestamp 1649977179
transform 1 0 61364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _529_
timestamp 1649977179
transform 1 0 60628 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _530__46
timestamp 1649977179
transform 1 0 27324 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _530_
timestamp 1649977179
transform 1 0 27140 0 1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _531__47
timestamp 1649977179
transform 1 0 63480 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _531_
timestamp 1649977179
transform 1 0 63204 0 1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _532__48
timestamp 1649977179
transform 1 0 32108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _532_
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _533__49
timestamp 1649977179
transform 1 0 38180 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _533_
timestamp 1649977179
transform 1 0 38088 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _534_
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _534__50
timestamp 1649977179
transform 1 0 36248 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _535__51
timestamp 1649977179
transform 1 0 42688 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _535_
timestamp 1649977179
transform 1 0 42596 0 -1 65280
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _536__52
timestamp 1649977179
transform 1 0 65596 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _536_
timestamp 1649977179
transform 1 0 65136 0 -1 62016
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _537__53
timestamp 1649977179
transform 1 0 43056 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _537_
timestamp 1649977179
transform 1 0 43424 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _538__54
timestamp 1649977179
transform 1 0 28152 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _538_
timestamp 1649977179
transform 1 0 28336 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _539__55
timestamp 1649977179
transform 1 0 30084 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _539_
timestamp 1649977179
transform 1 0 29716 0 -1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _540_
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _540__56
timestamp 1649977179
transform 1 0 54556 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _541__57
timestamp 1649977179
transform 1 0 51244 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _541_
timestamp 1649977179
transform 1 0 51152 0 1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _542__58
timestamp 1649977179
transform 1 0 26036 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _542_
timestamp 1649977179
transform 1 0 26036 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _543_
timestamp 1649977179
transform 1 0 43884 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _544__59
timestamp 1649977179
transform 1 0 55752 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _544_
timestamp 1649977179
transform 1 0 55660 0 1 64192
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _545__60
timestamp 1649977179
transform 1 0 46552 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _545_
timestamp 1649977179
transform 1 0 46460 0 1 62016
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _546__61
timestamp 1649977179
transform 1 0 67436 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _546_
timestamp 1649977179
transform 1 0 66240 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _547__62
timestamp 1649977179
transform 1 0 45356 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _547_
timestamp 1649977179
transform 1 0 45172 0 -1 51136
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _548_
timestamp 1649977179
transform 1 0 66240 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _548__63
timestamp 1649977179
transform 1 0 67436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _549__64
timestamp 1649977179
transform 1 0 67712 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _549_
timestamp 1649977179
transform 1 0 65780 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _550__65
timestamp 1649977179
transform 1 0 46552 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _550_
timestamp 1649977179
transform 1 0 46460 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _551__66
timestamp 1649977179
transform 1 0 51060 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _551_
timestamp 1649977179
transform 1 0 50968 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _552__67
timestamp 1649977179
transform 1 0 30084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _552_
timestamp 1649977179
transform 1 0 30084 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _553__68
timestamp 1649977179
transform 1 0 43884 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _553_
timestamp 1649977179
transform 1 0 43792 0 -1 66368
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _554_
timestamp 1649977179
transform 1 0 32108 0 -1 65280
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _554__69
timestamp 1649977179
transform 1 0 30728 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _555__70
timestamp 1649977179
transform 1 0 26220 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _555_
timestamp 1649977179
transform 1 0 26956 0 -1 59840
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _556__71
timestamp 1649977179
transform 1 0 37536 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _556_
timestamp 1649977179
transform 1 0 37444 0 -1 66368
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _557_
timestamp 1649977179
transform 1 0 27048 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _557__72
timestamp 1649977179
transform 1 0 27048 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _558__73
timestamp 1649977179
transform 1 0 10120 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _558_
timestamp 1649977179
transform 1 0 9200 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _559__74
timestamp 1649977179
transform 1 0 63388 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _559_
timestamp 1649977179
transform 1 0 63388 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _560__75
timestamp 1649977179
transform 1 0 43700 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _560_
timestamp 1649977179
transform 1 0 43608 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _561__76
timestamp 1649977179
transform 1 0 63296 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _561_
timestamp 1649977179
transform 1 0 63020 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _562__77
timestamp 1649977179
transform 1 0 7636 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _562_
timestamp 1649977179
transform 1 0 7544 0 -1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _563__78
timestamp 1649977179
transform 1 0 10488 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _563_
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _564_
timestamp 1649977179
transform 1 0 63112 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _564__79
timestamp 1649977179
transform 1 0 63112 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _565__80
timestamp 1649977179
transform 1 0 26772 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _565_
timestamp 1649977179
transform 1 0 26772 0 1 58752
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _566__81
timestamp 1649977179
transform 1 0 23000 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _566_
timestamp 1649977179
transform 1 0 23000 0 -1 60928
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _567_
timestamp 1649977179
transform 1 0 60904 0 1 67456
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _567__82
timestamp 1649977179
transform 1 0 61180 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _568_
timestamp 1649977179
transform 1 0 63020 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _568__83
timestamp 1649977179
transform 1 0 63020 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _569_
timestamp 1649977179
transform 1 0 8004 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _569__84
timestamp 1649977179
transform 1 0 8004 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _570__85
timestamp 1649977179
transform 1 0 50140 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _570_
timestamp 1649977179
transform 1 0 49680 0 -1 63104
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _571__86
timestamp 1649977179
transform 1 0 54096 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _571_
timestamp 1649977179
transform 1 0 54740 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _572__87
timestamp 1649977179
transform 1 0 38824 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _572_
timestamp 1649977179
transform 1 0 38824 0 -1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _573_
timestamp 1649977179
transform 1 0 52716 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _573__88
timestamp 1649977179
transform 1 0 52808 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _574__89
timestamp 1649977179
transform 1 0 53912 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _574_
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _575__90
timestamp 1649977179
transform 1 0 63664 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _575_
timestamp 1649977179
transform 1 0 63204 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _576__91
timestamp 1649977179
transform 1 0 4784 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _576_
timestamp 1649977179
transform 1 0 5060 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _577__92
timestamp 1649977179
transform 1 0 33580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _577_
timestamp 1649977179
transform 1 0 34224 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _578__93
timestamp 1649977179
transform 1 0 51428 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _578_
timestamp 1649977179
transform 1 0 51336 0 1 51136
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _579__94
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _579_
timestamp 1649977179
transform 1 0 19412 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _580__95
timestamp 1649977179
transform 1 0 26128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _580_
timestamp 1649977179
transform 1 0 26036 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _581__96
timestamp 1649977179
transform 1 0 24564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _581_
timestamp 1649977179
transform 1 0 24564 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _582__97
timestamp 1649977179
transform 1 0 67436 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _582_
timestamp 1649977179
transform 1 0 66240 0 1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _583__98
timestamp 1649977179
transform 1 0 56764 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _583_
timestamp 1649977179
transform 1 0 56212 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _584__99
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _584_
timestamp 1649977179
transform 1 0 34868 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _585_
timestamp 1649977179
transform 1 0 21988 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _585__100
timestamp 1649977179
transform 1 0 21988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _586_
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _586__101
timestamp 1649977179
transform 1 0 57684 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _587__102
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _587_
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _588__103
timestamp 1649977179
transform 1 0 4508 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _588_
timestamp 1649977179
transform 1 0 4508 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _589__104
timestamp 1649977179
transform 1 0 31372 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _589_
timestamp 1649977179
transform 1 0 32108 0 -1 63104
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _590__105
timestamp 1649977179
transform 1 0 31648 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _590_
timestamp 1649977179
transform 1 0 31648 0 1 64192
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _591__106
timestamp 1649977179
transform 1 0 59064 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _591_
timestamp 1649977179
transform 1 0 58972 0 -1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _592__107
timestamp 1649977179
transform 1 0 29992 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _592_
timestamp 1649977179
transform 1 0 32108 0 -1 64192
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _593__108
timestamp 1649977179
transform 1 0 54464 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _593_
timestamp 1649977179
transform 1 0 54464 0 -1 62016
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _594_
timestamp 1649977179
transform 1 0 65596 0 1 62016
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _594__109
timestamp 1649977179
transform 1 0 64860 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _595__110
timestamp 1649977179
transform 1 0 6256 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _595_
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _596__111
timestamp 1649977179
transform 1 0 57868 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _596_
timestamp 1649977179
transform 1 0 57592 0 1 63104
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _597_
timestamp 1649977179
transform 1 0 65320 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _597__112
timestamp 1649977179
transform 1 0 65596 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1649977179
transform 1 0 1380 0 -1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1649977179
transform 1 0 67344 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1649977179
transform 1 0 55476 0 -1 69632
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1649977179
transform 1 0 1380 0 -1 60928
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  repeater5
timestamp 1649977179
transform 1 0 32292 0 1 65280
box -38 -48 590 592
<< labels >>
flabel metal3 s 0 71348 800 71588 0 FreeSans 960 0 0 0 active
port 0 nsew signal input
flabel metal3 s 69200 22388 70000 22628 0 FreeSans 960 0 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 52154 0 52266 800 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 54730 0 54842 800 0 FreeSans 448 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 16090 0 16202 800 0 FreeSans 448 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal3 s 69200 11508 70000 11748 0 FreeSans 960 0 0 0 io_in[13]
port 5 nsew signal input
flabel metal3 s 69200 8788 70000 9028 0 FreeSans 960 0 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 25750 0 25862 800 0 FreeSans 448 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal3 s 0 10148 800 10388 0 FreeSans 960 0 0 0 io_in[16]
port 8 nsew signal input
flabel metal3 s 69200 36668 70000 36908 0 FreeSans 960 0 0 0 io_in[17]
port 9 nsew signal input
flabel metal3 s 69200 27148 70000 27388 0 FreeSans 960 0 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 57306 0 57418 800 0 FreeSans 448 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 21886 71200 21998 72000 0 FreeSans 448 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal3 s 69200 1988 70000 2228 0 FreeSans 960 0 0 0 io_in[20]
port 13 nsew signal input
flabel metal3 s 69200 52308 70000 52548 0 FreeSans 960 0 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 9006 71200 9118 72000 0 FreeSans 448 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 59238 71200 59350 72000 0 FreeSans 448 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal3 s 0 48228 800 48468 0 FreeSans 960 0 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 64390 71200 64502 72000 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 32834 71200 32946 72000 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 53442 0 53554 800 0 FreeSans 448 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal3 s 0 8788 800 9028 0 FreeSans 960 0 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 45714 0 45826 800 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 12870 71200 12982 72000 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 1278 71200 1390 72000 0 FreeSans 448 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 18022 71200 18134 72000 0 FreeSans 448 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal3 s 0 28508 800 28748 0 FreeSans 960 0 0 0 io_in[32]
port 26 nsew signal input
flabel metal3 s 69200 3348 70000 3588 0 FreeSans 960 0 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 37342 0 37454 800 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal3 s 69200 24428 70000 24668 0 FreeSans 960 0 0 0 io_in[35]
port 29 nsew signal input
flabel metal3 s 0 64548 800 64788 0 FreeSans 960 0 0 0 io_in[36]
port 30 nsew signal input
flabel metal3 s 69200 48228 70000 48468 0 FreeSans 960 0 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 59882 0 59994 800 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal3 s 0 57748 800 57988 0 FreeSans 960 0 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 23174 0 23286 800 0 FreeSans 448 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 30902 0 31014 800 0 FreeSans 448 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 58594 0 58706 800 0 FreeSans 448 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal3 s 0 14228 800 14468 0 FreeSans 960 0 0 0 io_in[8]
port 37 nsew signal input
flabel metal3 s 0 6068 800 6308 0 FreeSans 960 0 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 47002 0 47114 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal bidirectional
flabel metal2 s 50222 71200 50334 72000 0 FreeSans 448 90 0 0 io_oeb[10]
port 40 nsew signal bidirectional
flabel metal2 s 62458 0 62570 800 0 FreeSans 448 90 0 0 io_oeb[11]
port 41 nsew signal bidirectional
flabel metal2 s 52798 71200 52910 72000 0 FreeSans 448 90 0 0 io_oeb[12]
port 42 nsew signal bidirectional
flabel metal3 s 69200 43468 70000 43708 0 FreeSans 960 0 0 0 io_oeb[13]
port 43 nsew signal bidirectional
flabel metal3 s 69200 57748 70000 57988 0 FreeSans 960 0 0 0 io_oeb[14]
port 44 nsew signal bidirectional
flabel metal3 s 69200 42108 70000 42348 0 FreeSans 960 0 0 0 io_oeb[15]
port 45 nsew signal bidirectional
flabel metal3 s 0 23748 800 23988 0 FreeSans 960 0 0 0 io_oeb[16]
port 46 nsew signal bidirectional
flabel metal2 s 34766 0 34878 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal bidirectional
flabel metal2 s 63102 71200 63214 72000 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal bidirectional
flabel metal3 s 0 12868 800 13108 0 FreeSans 960 0 0 0 io_oeb[19]
port 49 nsew signal bidirectional
flabel metal3 s 69200 4708 70000 4948 0 FreeSans 960 0 0 0 io_oeb[1]
port 50 nsew signal bidirectional
flabel metal3 s 0 628 800 868 0 FreeSans 960 0 0 0 io_oeb[20]
port 51 nsew signal bidirectional
flabel metal2 s 19954 0 20066 800 0 FreeSans 448 90 0 0 io_oeb[21]
port 52 nsew signal bidirectional
flabel metal3 s 69200 65908 70000 66148 0 FreeSans 960 0 0 0 io_oeb[22]
port 53 nsew signal bidirectional
flabel metal2 s 56662 71200 56774 72000 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal bidirectional
flabel metal2 s 5786 0 5898 800 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal bidirectional
flabel metal2 s 22530 0 22642 800 0 FreeSans 448 90 0 0 io_oeb[25]
port 56 nsew signal bidirectional
flabel metal3 s 69200 40748 70000 40988 0 FreeSans 960 0 0 0 io_oeb[26]
port 57 nsew signal bidirectional
flabel metal2 s 45070 0 45182 800 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal bidirectional
flabel metal3 s 0 22388 800 22628 0 FreeSans 960 0 0 0 io_oeb[28]
port 59 nsew signal bidirectional
flabel metal2 s 31546 71200 31658 72000 0 FreeSans 448 90 0 0 io_oeb[29]
port 60 nsew signal bidirectional
flabel metal3 s 0 52308 800 52548 0 FreeSans 960 0 0 0 io_oeb[2]
port 61 nsew signal bidirectional
flabel metal2 s 5142 71200 5254 72000 0 FreeSans 448 90 0 0 io_oeb[30]
port 62 nsew signal bidirectional
flabel metal2 s 68254 71200 68366 72000 0 FreeSans 448 90 0 0 io_oeb[31]
port 63 nsew signal bidirectional
flabel metal2 s 39274 71200 39386 72000 0 FreeSans 448 90 0 0 io_oeb[32]
port 64 nsew signal bidirectional
flabel metal3 s 69200 61828 70000 62068 0 FreeSans 960 0 0 0 io_oeb[33]
port 65 nsew signal bidirectional
flabel metal3 s 69200 63188 70000 63428 0 FreeSans 960 0 0 0 io_oeb[34]
port 66 nsew signal bidirectional
flabel metal3 s 0 35308 800 35548 0 FreeSans 960 0 0 0 io_oeb[35]
port 67 nsew signal bidirectional
flabel metal2 s 57950 71200 58062 72000 0 FreeSans 448 90 0 0 io_oeb[36]
port 68 nsew signal bidirectional
flabel metal3 s 69200 46188 70000 46428 0 FreeSans 960 0 0 0 io_oeb[37]
port 69 nsew signal bidirectional
flabel metal2 s 11582 71200 11694 72000 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal bidirectional
flabel metal3 s 69200 21028 70000 21268 0 FreeSans 960 0 0 0 io_oeb[4]
port 71 nsew signal bidirectional
flabel metal3 s 0 59108 800 59348 0 FreeSans 960 0 0 0 io_oeb[5]
port 72 nsew signal bidirectional
flabel metal2 s 6430 71200 6542 72000 0 FreeSans 448 90 0 0 io_oeb[6]
port 73 nsew signal bidirectional
flabel metal3 s 69200 67268 70000 67508 0 FreeSans 960 0 0 0 io_oeb[7]
port 74 nsew signal bidirectional
flabel metal3 s 69200 35308 70000 35548 0 FreeSans 960 0 0 0 io_oeb[8]
port 75 nsew signal bidirectional
flabel metal3 s 0 29868 800 30108 0 FreeSans 960 0 0 0 io_oeb[9]
port 76 nsew signal bidirectional
flabel metal3 s 0 67268 800 67508 0 FreeSans 960 0 0 0 io_out[0]
port 77 nsew signal bidirectional
flabel metal3 s 0 1988 800 2228 0 FreeSans 960 0 0 0 io_out[10]
port 78 nsew signal bidirectional
flabel metal2 s 38630 0 38742 800 0 FreeSans 448 90 0 0 io_out[11]
port 79 nsew signal bidirectional
flabel metal3 s 0 31228 800 31468 0 FreeSans 960 0 0 0 io_out[12]
port 80 nsew signal bidirectional
flabel metal2 s 43138 71200 43250 72000 0 FreeSans 448 90 0 0 io_out[13]
port 81 nsew signal bidirectional
flabel metal2 s 69542 71200 69654 72000 0 FreeSans 448 90 0 0 io_out[14]
port 82 nsew signal bidirectional
flabel metal3 s 0 47548 800 47788 0 FreeSans 960 0 0 0 io_out[15]
port 83 nsew signal bidirectional
flabel metal2 s 7074 0 7186 800 0 FreeSans 448 90 0 0 io_out[16]
port 84 nsew signal bidirectional
flabel metal2 s 25106 71200 25218 72000 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal bidirectional
flabel metal3 s 69200 16948 70000 17188 0 FreeSans 960 0 0 0 io_out[18]
port 86 nsew signal bidirectional
flabel metal2 s 60526 71200 60638 72000 0 FreeSans 448 90 0 0 io_out[19]
port 87 nsew signal bidirectional
flabel metal3 s 0 3348 800 3588 0 FreeSans 960 0 0 0 io_out[1]
port 88 nsew signal bidirectional
flabel metal3 s 0 25788 800 26028 0 FreeSans 960 0 0 0 io_out[20]
port 89 nsew signal bidirectional
flabel metal2 s 61170 0 61282 800 0 FreeSans 448 90 0 0 io_out[21]
port 90 nsew signal bidirectional
flabel metal2 s 66966 71200 67078 72000 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal bidirectional
flabel metal2 s 47002 71200 47114 72000 0 FreeSans 448 90 0 0 io_out[23]
port 92 nsew signal bidirectional
flabel metal3 s 69200 44828 70000 45068 0 FreeSans 960 0 0 0 io_out[24]
port 93 nsew signal bidirectional
flabel metal3 s 0 53668 800 53908 0 FreeSans 960 0 0 0 io_out[25]
port 94 nsew signal bidirectional
flabel metal2 s 69542 0 69654 800 0 FreeSans 448 90 0 0 io_out[26]
port 95 nsew signal bidirectional
flabel metal3 s 69200 31228 70000 31468 0 FreeSans 960 0 0 0 io_out[27]
port 96 nsew signal bidirectional
flabel metal2 s 41850 71200 41962 72000 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal bidirectional
flabel metal2 s 51510 71200 51622 72000 0 FreeSans 448 90 0 0 io_out[29]
port 98 nsew signal bidirectional
flabel metal3 s 69200 23068 70000 23308 0 FreeSans 960 0 0 0 io_out[2]
port 99 nsew signal bidirectional
flabel metal3 s 0 4708 800 4948 0 FreeSans 960 0 0 0 io_out[30]
port 100 nsew signal bidirectional
flabel metal2 s 45714 71200 45826 72000 0 FreeSans 448 90 0 0 io_out[31]
port 101 nsew signal bidirectional
flabel metal2 s 16734 71200 16846 72000 0 FreeSans 448 90 0 0 io_out[32]
port 102 nsew signal bidirectional
flabel metal2 s 27682 71200 27794 72000 0 FreeSans 448 90 0 0 io_out[33]
port 103 nsew signal bidirectional
flabel metal2 s 37986 71200 38098 72000 0 FreeSans 448 90 0 0 io_out[34]
port 104 nsew signal bidirectional
flabel metal2 s 68898 0 69010 800 0 FreeSans 448 90 0 0 io_out[35]
port 105 nsew signal bidirectional
flabel metal3 s 0 15588 800 15828 0 FreeSans 960 0 0 0 io_out[36]
port 106 nsew signal bidirectional
flabel metal3 s 69200 6068 70000 6308 0 FreeSans 960 0 0 0 io_out[37]
port 107 nsew signal bidirectional
flabel metal2 s 10938 0 11050 800 0 FreeSans 448 90 0 0 io_out[3]
port 108 nsew signal bidirectional
flabel metal3 s 0 39388 800 39628 0 FreeSans 960 0 0 0 io_out[4]
port 109 nsew signal bidirectional
flabel metal2 s 36698 71200 36810 72000 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal bidirectional
flabel metal3 s 69200 32588 70000 32828 0 FreeSans 960 0 0 0 io_out[6]
port 111 nsew signal bidirectional
flabel metal3 s 69200 14228 70000 14468 0 FreeSans 960 0 0 0 io_out[7]
port 112 nsew signal bidirectional
flabel metal3 s 0 68628 800 68868 0 FreeSans 960 0 0 0 io_out[8]
port 113 nsew signal bidirectional
flabel metal3 s 69200 60468 70000 60708 0 FreeSans 960 0 0 0 io_out[9]
port 114 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 69680 0 FreeSans 1920 90 0 0 vccd1
port 115 nsew power bidirectional
flabel metal4 s 34928 2128 35248 69680 0 FreeSans 1920 90 0 0 vccd1
port 115 nsew power bidirectional
flabel metal4 s 65648 2128 65968 69680 0 FreeSans 1920 90 0 0 vccd1
port 115 nsew power bidirectional
flabel metal4 s 19568 2128 19888 69680 0 FreeSans 1920 90 0 0 vssd1
port 116 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 69680 0 FreeSans 1920 90 0 0 vssd1
port 116 nsew ground bidirectional
flabel metal2 s 23174 71200 23286 72000 0 FreeSans 448 90 0 0 wb_clk_i
port 117 nsew signal input
flabel metal3 s 69200 69988 70000 70228 0 FreeSans 960 0 0 0 wb_rst_i
port 118 nsew signal input
flabel metal3 s 0 50948 800 51188 0 FreeSans 960 0 0 0 wbs_ack_o
port 119 nsew signal bidirectional
flabel metal3 s 69200 47548 70000 47788 0 FreeSans 960 0 0 0 wbs_adr_i[0]
port 120 nsew signal input
flabel metal3 s 69200 59108 70000 59348 0 FreeSans 960 0 0 0 wbs_adr_i[10]
port 121 nsew signal input
flabel metal3 s 0 42108 800 42348 0 FreeSans 960 0 0 0 wbs_adr_i[11]
port 122 nsew signal input
flabel metal2 s 3210 0 3322 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 123 nsew signal input
flabel metal2 s 27038 0 27150 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 124 nsew signal input
flabel metal3 s 69200 18308 70000 18548 0 FreeSans 960 0 0 0 wbs_adr_i[14]
port 125 nsew signal input
flabel metal2 s 35410 71200 35522 72000 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 126 nsew signal input
flabel metal2 s 32190 0 32302 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 127 nsew signal input
flabel metal3 s 69200 12868 70000 13108 0 FreeSans 960 0 0 0 wbs_adr_i[17]
port 128 nsew signal input
flabel metal2 s 67610 0 67722 800 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 129 nsew signal input
flabel metal3 s 0 63188 800 63428 0 FreeSans 960 0 0 0 wbs_adr_i[19]
port 130 nsew signal input
flabel metal3 s 0 46188 800 46428 0 FreeSans 960 0 0 0 wbs_adr_i[1]
port 131 nsew signal input
flabel metal3 s 69200 39388 70000 39628 0 FreeSans 960 0 0 0 wbs_adr_i[20]
port 132 nsew signal input
flabel metal3 s 0 56388 800 56628 0 FreeSans 960 0 0 0 wbs_adr_i[21]
port 133 nsew signal input
flabel metal3 s 0 24428 800 24668 0 FreeSans 960 0 0 0 wbs_adr_i[22]
port 134 nsew signal input
flabel metal2 s 65034 0 65146 800 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 135 nsew signal input
flabel metal2 s 20598 71200 20710 72000 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 136 nsew signal input
flabel metal2 s 28326 0 28438 800 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 137 nsew signal input
flabel metal3 s 0 33948 800 34188 0 FreeSans 960 0 0 0 wbs_adr_i[26]
port 138 nsew signal input
flabel metal3 s 0 44828 800 45068 0 FreeSans 960 0 0 0 wbs_adr_i[27]
port 139 nsew signal input
flabel metal3 s 0 21028 800 21268 0 FreeSans 960 0 0 0 wbs_adr_i[28]
port 140 nsew signal input
flabel metal2 s 19310 71200 19422 72000 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 141 nsew signal input
flabel metal2 s 21242 0 21354 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 142 nsew signal input
flabel metal2 s 7718 71200 7830 72000 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 143 nsew signal input
flabel metal3 s 69200 7428 70000 7668 0 FreeSans 960 0 0 0 wbs_adr_i[31]
port 144 nsew signal input
flabel metal2 s 42494 0 42606 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 145 nsew signal input
flabel metal3 s 69200 56388 70000 56628 0 FreeSans 960 0 0 0 wbs_adr_i[4]
port 146 nsew signal input
flabel metal3 s 0 7428 800 7668 0 FreeSans 960 0 0 0 wbs_adr_i[5]
port 147 nsew signal input
flabel metal2 s 17378 0 17490 800 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 148 nsew signal input
flabel metal2 s 14158 71200 14270 72000 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 149 nsew signal input
flabel metal2 s 56018 0 56130 800 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 150 nsew signal input
flabel metal3 s 0 43468 800 43708 0 FreeSans 960 0 0 0 wbs_adr_i[9]
port 151 nsew signal input
flabel metal2 s 55374 71200 55486 72000 0 FreeSans 448 90 0 0 wbs_cyc_i
port 152 nsew signal input
flabel metal2 s 634 71200 746 72000 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 153 nsew signal input
flabel metal2 s 15446 71200 15558 72000 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 154 nsew signal input
flabel metal2 s 26394 71200 26506 72000 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 155 nsew signal input
flabel metal2 s 23818 71200 23930 72000 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 156 nsew signal input
flabel metal2 s 1922 0 2034 800 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 157 nsew signal input
flabel metal2 s 12226 0 12338 800 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 158 nsew signal input
flabel metal3 s 0 19668 800 19908 0 FreeSans 960 0 0 0 wbs_dat_i[15]
port 159 nsew signal input
flabel metal2 s 33478 0 33590 800 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 160 nsew signal input
flabel metal3 s 69200 68628 70000 68868 0 FreeSans 960 0 0 0 wbs_dat_i[17]
port 161 nsew signal input
flabel metal2 s 2566 71200 2678 72000 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 162 nsew signal input
flabel metal2 s 34122 71200 34234 72000 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 163 nsew signal input
flabel metal2 s 8362 0 8474 800 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 164 nsew signal input
flabel metal3 s 69200 25788 70000 26028 0 FreeSans 960 0 0 0 wbs_dat_i[20]
port 165 nsew signal input
flabel metal3 s 69200 53668 70000 53908 0 FreeSans 960 0 0 0 wbs_dat_i[21]
port 166 nsew signal input
flabel metal3 s 0 32588 800 32828 0 FreeSans 960 0 0 0 wbs_dat_i[22]
port 167 nsew signal input
flabel metal3 s 69200 38028 70000 38268 0 FreeSans 960 0 0 0 wbs_dat_i[23]
port 168 nsew signal input
flabel metal3 s 0 61828 800 62068 0 FreeSans 960 0 0 0 wbs_dat_i[24]
port 169 nsew signal input
flabel metal3 s 0 11508 800 11748 0 FreeSans 960 0 0 0 wbs_dat_i[25]
port 170 nsew signal input
flabel metal3 s 69200 64548 70000 64788 0 FreeSans 960 0 0 0 wbs_dat_i[26]
port 171 nsew signal input
flabel metal2 s 40562 71200 40674 72000 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 172 nsew signal input
flabel metal2 s 18666 0 18778 800 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 173 nsew signal input
flabel metal3 s 69200 28508 70000 28748 0 FreeSans 960 0 0 0 wbs_dat_i[29]
port 174 nsew signal input
flabel metal2 s 49578 0 49690 800 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 175 nsew signal input
flabel metal3 s 69200 10148 70000 10388 0 FreeSans 960 0 0 0 wbs_dat_i[30]
port 176 nsew signal input
flabel metal3 s 0 65908 800 66148 0 FreeSans 960 0 0 0 wbs_dat_i[31]
port 177 nsew signal input
flabel metal2 s 63746 0 63858 800 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 178 nsew signal input
flabel metal2 s 9650 0 9762 800 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 179 nsew signal input
flabel metal2 s 29614 0 29726 800 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 180 nsew signal input
flabel metal3 s 69200 19668 70000 19908 0 FreeSans 960 0 0 0 wbs_dat_i[6]
port 181 nsew signal input
flabel metal3 s 69200 71348 70000 71588 0 FreeSans 960 0 0 0 wbs_dat_i[7]
port 182 nsew signal input
flabel metal3 s 0 18308 800 18548 0 FreeSans 960 0 0 0 wbs_dat_i[8]
port 183 nsew signal input
flabel metal2 s 66322 0 66434 800 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 184 nsew signal input
flabel metal3 s 0 27148 800 27388 0 FreeSans 960 0 0 0 wbs_dat_o[0]
port 185 nsew signal bidirectional
flabel metal3 s 69200 29868 70000 30108 0 FreeSans 960 0 0 0 wbs_dat_o[10]
port 186 nsew signal bidirectional
flabel metal2 s 634 0 746 800 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 187 nsew signal bidirectional
flabel metal3 s 69200 55028 70000 55268 0 FreeSans 960 0 0 0 wbs_dat_o[12]
port 188 nsew signal bidirectional
flabel metal2 s 65678 71200 65790 72000 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 189 nsew signal bidirectional
flabel metal3 s 69200 628 70000 868 0 FreeSans 960 0 0 0 wbs_dat_o[14]
port 190 nsew signal bidirectional
flabel metal2 s 61814 71200 61926 72000 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 191 nsew signal bidirectional
flabel metal3 s 0 38028 800 38268 0 FreeSans 960 0 0 0 wbs_dat_o[16]
port 192 nsew signal bidirectional
flabel metal3 s 0 40748 800 40988 0 FreeSans 960 0 0 0 wbs_dat_o[17]
port 193 nsew signal bidirectional
flabel metal2 s 43782 0 43894 800 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 194 nsew signal bidirectional
flabel metal2 s -10 0 102 800 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 195 nsew signal bidirectional
flabel metal2 s 50866 0 50978 800 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 196 nsew signal bidirectional
flabel metal3 s 0 49588 800 49828 0 FreeSans 960 0 0 0 wbs_dat_o[20]
port 197 nsew signal bidirectional
flabel metal2 s 3854 71200 3966 72000 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 198 nsew signal bidirectional
flabel metal2 s 30258 71200 30370 72000 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 199 nsew signal bidirectional
flabel metal3 s 0 36668 800 36908 0 FreeSans 960 0 0 0 wbs_dat_o[23]
port 200 nsew signal bidirectional
flabel metal2 s 13514 0 13626 800 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 201 nsew signal bidirectional
flabel metal2 s 4498 0 4610 800 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 202 nsew signal bidirectional
flabel metal2 s 44426 71200 44538 72000 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 203 nsew signal bidirectional
flabel metal2 s 28970 71200 29082 72000 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 204 nsew signal bidirectional
flabel metal2 s 36054 0 36166 800 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 205 nsew signal bidirectional
flabel metal2 s 54086 71200 54198 72000 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 206 nsew signal bidirectional
flabel metal3 s 69200 15588 70000 15828 0 FreeSans 960 0 0 0 wbs_dat_o[2]
port 207 nsew signal bidirectional
flabel metal3 s 0 55028 800 55268 0 FreeSans 960 0 0 0 wbs_dat_o[30]
port 208 nsew signal bidirectional
flabel metal3 s 69200 50948 70000 51188 0 FreeSans 960 0 0 0 wbs_dat_o[31]
port 209 nsew signal bidirectional
flabel metal2 s 14802 0 14914 800 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 210 nsew signal bidirectional
flabel metal2 s 24462 0 24574 800 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 211 nsew signal bidirectional
flabel metal2 s 39918 0 40030 800 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 212 nsew signal bidirectional
flabel metal3 s 69200 49588 70000 49828 0 FreeSans 960 0 0 0 wbs_dat_o[6]
port 213 nsew signal bidirectional
flabel metal2 s 41206 0 41318 800 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 214 nsew signal bidirectional
flabel metal2 s 48934 71200 49046 72000 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 215 nsew signal bidirectional
flabel metal2 s 47646 71200 47758 72000 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 216 nsew signal bidirectional
flabel metal3 s 0 69988 800 70228 0 FreeSans 960 0 0 0 wbs_sel_i[0]
port 217 nsew signal input
flabel metal2 s 10294 71200 10406 72000 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 218 nsew signal input
flabel metal2 s 48290 0 48402 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 219 nsew signal input
flabel metal3 s 0 16948 800 17188 0 FreeSans 960 0 0 0 wbs_sel_i[3]
port 220 nsew signal input
flabel metal3 s 0 60468 800 60708 0 FreeSans 960 0 0 0 wbs_stb_i
port 221 nsew signal input
flabel metal3 s 69200 33948 70000 34188 0 FreeSans 960 0 0 0 wbs_we_i
port 222 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 72000
<< end >>
