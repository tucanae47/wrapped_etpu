VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_etpu
  CLASS BLOCK ;
  FOREIGN wrapped_etpu ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 360.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.340 4.000 354.540 ;
    END
  END active
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 348.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 348.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 348.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 348.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 348.400 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 349.940 350.000 351.140 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 0.000 206.590 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 0.000 103.550 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.740 4.000 204.940 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 356.000 213.030 360.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.390 356.000 328.950 360.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.110 356.000 251.670 360.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.940 4.000 28.140 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 356.000 174.390 360.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.950 0.000 322.510 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 200.340 350.000 201.540 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 0.000 77.790 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.740 4.000 272.940 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.230 356.000 238.790 360.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.070 0.000 309.630 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 0.000 142.190 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 309.140 350.000 310.340 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.940 4.000 300.140 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 118.740 350.000 119.940 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 295.540 350.000 296.740 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.750 356.000 290.310 360.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 77.940 350.000 79.140 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 336.340 350.000 337.540 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.740 4.000 68.940 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.340 4.000 150.540 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 64.340 350.000 65.540 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.140 4.000 191.340 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.540 4.000 245.740 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 356.000 97.110 360.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 356.000 187.270 360.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.510 356.000 316.070 360.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 0.000 39.150 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 268.340 350.000 269.540 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.940 4.000 232.140 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 23.540 350.000 24.740 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.430 0.000 270.990 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 159.540 350.000 160.740 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 132.340 350.000 133.540 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 356.000 109.990 360.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 356.000 122.870 360.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 281.940 350.000 283.140 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.140 4.000 55.340 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 0.000 90.670 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 50.740 350.000 51.940 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 9.940 350.000 11.140 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 186.740 350.000 187.940 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.140 4.000 259.340 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.190 0.000 296.750 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 356.000 135.750 360.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 322.740 350.000 323.940 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.710 0.000 348.270 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.950 356.000 161.510 360.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 0.000 129.310 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 91.540 350.000 92.740 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 227.540 350.000 228.740 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.540 4.000 177.740 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 356.000 200.150 360.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.390 0.000 167.950 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 356.000 84.230 360.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.140 4.000 327.340 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 0.000 232.350 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 0.000 26.270 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.940 4.000 164.140 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.830 0.000 335.390 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 105.140 350.000 106.340 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.550 0.000 258.110 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.340 4.000 286.540 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.340 4.000 218.540 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.340 4.000 82.540 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 145.940 350.000 147.140 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 241.140 350.000 242.340 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 0.000 283.870 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 254.740 350.000 255.940 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 356.000 32.710 360.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030 356.000 45.590 360.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 0.000 180.830 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 0.000 219.470 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 356.000 58.470 360.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 356.000 148.630 360.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.940 4.000 96.140 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.740 4.000 340.940 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 0.000 52.030 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 0.000 13.390 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.630 356.000 303.190 360.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.350 356.000 225.910 360.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.510 0.000 155.070 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 356.000 341.830 360.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 37.140 350.000 38.340 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 356.000 6.950 360.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.740 4.000 136.940 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 0.000 64.910 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 0.000 116.430 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.140 4.000 123.340 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 213.940 350.000 215.140 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 0.000 193.710 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.870 356.000 277.430 360.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 356.000 264.550 360.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.270 356.000 19.830 360.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 356.000 71.350 360.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 0.000 245.230 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.540 4.000 109.740 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.540 4.000 313.740 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 173.140 350.000 174.340 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 348.245 ;
      LAYER met1 ;
        RECT 0.070 10.640 344.080 348.400 ;
      LAYER met2 ;
        RECT 0.100 355.720 6.110 356.000 ;
        RECT 7.230 355.720 18.990 356.000 ;
        RECT 20.110 355.720 31.870 356.000 ;
        RECT 32.990 355.720 44.750 356.000 ;
        RECT 45.870 355.720 57.630 356.000 ;
        RECT 58.750 355.720 70.510 356.000 ;
        RECT 71.630 355.720 83.390 356.000 ;
        RECT 84.510 355.720 96.270 356.000 ;
        RECT 97.390 355.720 109.150 356.000 ;
        RECT 110.270 355.720 122.030 356.000 ;
        RECT 123.150 355.720 134.910 356.000 ;
        RECT 136.030 355.720 147.790 356.000 ;
        RECT 148.910 355.720 160.670 356.000 ;
        RECT 161.790 355.720 173.550 356.000 ;
        RECT 174.670 355.720 186.430 356.000 ;
        RECT 187.550 355.720 199.310 356.000 ;
        RECT 200.430 355.720 212.190 356.000 ;
        RECT 213.310 355.720 225.070 356.000 ;
        RECT 226.190 355.720 237.950 356.000 ;
        RECT 239.070 355.720 250.830 356.000 ;
        RECT 251.950 355.720 263.710 356.000 ;
        RECT 264.830 355.720 276.590 356.000 ;
        RECT 277.710 355.720 289.470 356.000 ;
        RECT 290.590 355.720 302.350 356.000 ;
        RECT 303.470 355.720 315.230 356.000 ;
        RECT 316.350 355.720 328.110 356.000 ;
        RECT 329.230 355.720 340.990 356.000 ;
        RECT 0.100 4.280 341.680 355.720 ;
        RECT 0.790 3.670 12.550 4.280 ;
        RECT 13.670 3.670 25.430 4.280 ;
        RECT 26.550 3.670 38.310 4.280 ;
        RECT 39.430 3.670 51.190 4.280 ;
        RECT 52.310 3.670 64.070 4.280 ;
        RECT 65.190 3.670 76.950 4.280 ;
        RECT 78.070 3.670 89.830 4.280 ;
        RECT 90.950 3.670 102.710 4.280 ;
        RECT 103.830 3.670 115.590 4.280 ;
        RECT 116.710 3.670 128.470 4.280 ;
        RECT 129.590 3.670 141.350 4.280 ;
        RECT 142.470 3.670 154.230 4.280 ;
        RECT 155.350 3.670 167.110 4.280 ;
        RECT 168.230 3.670 179.990 4.280 ;
        RECT 181.110 3.670 192.870 4.280 ;
        RECT 193.990 3.670 205.750 4.280 ;
        RECT 206.870 3.670 218.630 4.280 ;
        RECT 219.750 3.670 231.510 4.280 ;
        RECT 232.630 3.670 244.390 4.280 ;
        RECT 245.510 3.670 257.270 4.280 ;
        RECT 258.390 3.670 270.150 4.280 ;
        RECT 271.270 3.670 283.030 4.280 ;
        RECT 284.150 3.670 295.910 4.280 ;
        RECT 297.030 3.670 308.790 4.280 ;
        RECT 309.910 3.670 321.670 4.280 ;
        RECT 322.790 3.670 334.550 4.280 ;
        RECT 335.670 3.670 341.680 4.280 ;
      LAYER met3 ;
        RECT 4.400 352.940 346.000 354.105 ;
        RECT 4.000 351.540 346.000 352.940 ;
        RECT 4.000 349.540 345.600 351.540 ;
        RECT 4.000 341.340 346.000 349.540 ;
        RECT 4.400 339.340 346.000 341.340 ;
        RECT 4.000 337.940 346.000 339.340 ;
        RECT 4.000 335.940 345.600 337.940 ;
        RECT 4.000 327.740 346.000 335.940 ;
        RECT 4.400 325.740 346.000 327.740 ;
        RECT 4.000 324.340 346.000 325.740 ;
        RECT 4.000 322.340 345.600 324.340 ;
        RECT 4.000 314.140 346.000 322.340 ;
        RECT 4.400 312.140 346.000 314.140 ;
        RECT 4.000 310.740 346.000 312.140 ;
        RECT 4.000 308.740 345.600 310.740 ;
        RECT 4.000 300.540 346.000 308.740 ;
        RECT 4.400 298.540 346.000 300.540 ;
        RECT 4.000 297.140 346.000 298.540 ;
        RECT 4.000 295.140 345.600 297.140 ;
        RECT 4.000 286.940 346.000 295.140 ;
        RECT 4.400 284.940 346.000 286.940 ;
        RECT 4.000 283.540 346.000 284.940 ;
        RECT 4.000 281.540 345.600 283.540 ;
        RECT 4.000 273.340 346.000 281.540 ;
        RECT 4.400 271.340 346.000 273.340 ;
        RECT 4.000 269.940 346.000 271.340 ;
        RECT 4.000 267.940 345.600 269.940 ;
        RECT 4.000 259.740 346.000 267.940 ;
        RECT 4.400 257.740 346.000 259.740 ;
        RECT 4.000 256.340 346.000 257.740 ;
        RECT 4.000 254.340 345.600 256.340 ;
        RECT 4.000 246.140 346.000 254.340 ;
        RECT 4.400 244.140 346.000 246.140 ;
        RECT 4.000 242.740 346.000 244.140 ;
        RECT 4.000 240.740 345.600 242.740 ;
        RECT 4.000 232.540 346.000 240.740 ;
        RECT 4.400 230.540 346.000 232.540 ;
        RECT 4.000 229.140 346.000 230.540 ;
        RECT 4.000 227.140 345.600 229.140 ;
        RECT 4.000 218.940 346.000 227.140 ;
        RECT 4.400 216.940 346.000 218.940 ;
        RECT 4.000 215.540 346.000 216.940 ;
        RECT 4.000 213.540 345.600 215.540 ;
        RECT 4.000 205.340 346.000 213.540 ;
        RECT 4.400 203.340 346.000 205.340 ;
        RECT 4.000 201.940 346.000 203.340 ;
        RECT 4.000 199.940 345.600 201.940 ;
        RECT 4.000 191.740 346.000 199.940 ;
        RECT 4.400 189.740 346.000 191.740 ;
        RECT 4.000 188.340 346.000 189.740 ;
        RECT 4.000 186.340 345.600 188.340 ;
        RECT 4.000 178.140 346.000 186.340 ;
        RECT 4.400 176.140 346.000 178.140 ;
        RECT 4.000 174.740 346.000 176.140 ;
        RECT 4.000 172.740 345.600 174.740 ;
        RECT 4.000 164.540 346.000 172.740 ;
        RECT 4.400 162.540 346.000 164.540 ;
        RECT 4.000 161.140 346.000 162.540 ;
        RECT 4.000 159.140 345.600 161.140 ;
        RECT 4.000 150.940 346.000 159.140 ;
        RECT 4.400 148.940 346.000 150.940 ;
        RECT 4.000 147.540 346.000 148.940 ;
        RECT 4.000 145.540 345.600 147.540 ;
        RECT 4.000 137.340 346.000 145.540 ;
        RECT 4.400 135.340 346.000 137.340 ;
        RECT 4.000 133.940 346.000 135.340 ;
        RECT 4.000 131.940 345.600 133.940 ;
        RECT 4.000 123.740 346.000 131.940 ;
        RECT 4.400 121.740 346.000 123.740 ;
        RECT 4.000 120.340 346.000 121.740 ;
        RECT 4.000 118.340 345.600 120.340 ;
        RECT 4.000 110.140 346.000 118.340 ;
        RECT 4.400 108.140 346.000 110.140 ;
        RECT 4.000 106.740 346.000 108.140 ;
        RECT 4.000 104.740 345.600 106.740 ;
        RECT 4.000 96.540 346.000 104.740 ;
        RECT 4.400 94.540 346.000 96.540 ;
        RECT 4.000 93.140 346.000 94.540 ;
        RECT 4.000 91.140 345.600 93.140 ;
        RECT 4.000 82.940 346.000 91.140 ;
        RECT 4.400 80.940 346.000 82.940 ;
        RECT 4.000 79.540 346.000 80.940 ;
        RECT 4.000 77.540 345.600 79.540 ;
        RECT 4.000 69.340 346.000 77.540 ;
        RECT 4.400 67.340 346.000 69.340 ;
        RECT 4.000 65.940 346.000 67.340 ;
        RECT 4.000 63.940 345.600 65.940 ;
        RECT 4.000 55.740 346.000 63.940 ;
        RECT 4.400 53.740 346.000 55.740 ;
        RECT 4.000 52.340 346.000 53.740 ;
        RECT 4.000 50.340 345.600 52.340 ;
        RECT 4.000 42.140 346.000 50.340 ;
        RECT 4.400 40.140 346.000 42.140 ;
        RECT 4.000 38.740 346.000 40.140 ;
        RECT 4.000 36.740 345.600 38.740 ;
        RECT 4.000 28.540 346.000 36.740 ;
        RECT 4.400 26.540 346.000 28.540 ;
        RECT 4.000 25.140 346.000 26.540 ;
        RECT 4.000 23.140 345.600 25.140 ;
        RECT 4.000 14.940 346.000 23.140 ;
        RECT 4.400 12.940 346.000 14.940 ;
        RECT 4.000 11.540 346.000 12.940 ;
        RECT 4.000 10.715 345.600 11.540 ;
  END
END wrapped_etpu
END LIBRARY

