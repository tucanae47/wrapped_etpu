magic
tech sky130A
magscale 1 2
timestamp 1654694705
<< viali >>
rect 1409 66113 1443 66147
rect 1593 66045 1627 66079
rect 19809 64413 19843 64447
rect 21281 64005 21315 64039
rect 19441 63937 19475 63971
rect 19625 63869 19659 63903
rect 18981 63733 19015 63767
rect 19349 63393 19383 63427
rect 19809 63393 19843 63427
rect 43361 63325 43395 63359
rect 44005 63325 44039 63359
rect 19533 63257 19567 63291
rect 43453 63189 43487 63223
rect 19533 62985 19567 63019
rect 20177 62985 20211 63019
rect 43821 62917 43855 62951
rect 19625 62849 19659 62883
rect 20269 62849 20303 62883
rect 43637 62849 43671 62883
rect 45477 62781 45511 62815
rect 32781 62237 32815 62271
rect 37105 62237 37139 62271
rect 30941 62169 30975 62203
rect 32597 62169 32631 62203
rect 32229 61897 32263 61931
rect 32321 61761 32355 61795
rect 36553 61761 36587 61795
rect 37289 61761 37323 61795
rect 31217 61693 31251 61727
rect 36645 61693 36679 61727
rect 37473 61693 37507 61727
rect 37749 61693 37783 61727
rect 45937 61557 45971 61591
rect 54769 61557 54803 61591
rect 45845 61217 45879 61251
rect 46305 61217 46339 61251
rect 55321 61217 55355 61251
rect 54125 61149 54159 61183
rect 46029 61081 46063 61115
rect 54217 61081 54251 61115
rect 55505 61081 55539 61115
rect 57161 61081 57195 61115
rect 46029 60809 46063 60843
rect 45937 60673 45971 60707
rect 26525 60061 26559 60095
rect 35633 60061 35667 60095
rect 55321 60061 55355 60095
rect 54309 59653 54343 59687
rect 55045 59653 55079 59687
rect 56701 59653 56735 59687
rect 26249 59585 26283 59619
rect 26985 59585 27019 59619
rect 54217 59585 54251 59619
rect 54861 59585 54895 59619
rect 26341 59517 26375 59551
rect 27169 59517 27203 59551
rect 27445 59517 27479 59551
rect 35541 59041 35575 59075
rect 37197 59041 37231 59075
rect 35725 58905 35759 58939
rect 35725 58633 35759 58667
rect 66177 58565 66211 58599
rect 35633 58497 35667 58531
rect 37473 58497 37507 58531
rect 64337 58429 64371 58463
rect 64521 58429 64555 58463
rect 36553 58361 36587 58395
rect 37381 58293 37415 58327
rect 64705 58089 64739 58123
rect 65625 58089 65659 58123
rect 37933 57953 37967 57987
rect 34713 57885 34747 57919
rect 36277 57885 36311 57919
rect 38117 57885 38151 57919
rect 63509 57885 63543 57919
rect 63969 57885 64003 57919
rect 64613 57885 64647 57919
rect 64061 57749 64095 57783
rect 64245 57477 64279 57511
rect 65901 57477 65935 57511
rect 34253 57409 34287 57443
rect 64061 57409 64095 57443
rect 34437 57341 34471 57375
rect 35817 57341 35851 57375
rect 34805 57001 34839 57035
rect 34897 56797 34931 56831
rect 49249 56797 49283 56831
rect 64061 56797 64095 56831
rect 49249 56321 49283 56355
rect 63969 56321 64003 56355
rect 32965 56253 32999 56287
rect 33149 56253 33183 56287
rect 33425 56253 33459 56287
rect 49433 56253 49467 56287
rect 51089 56253 51123 56287
rect 64153 56253 64187 56287
rect 64429 56253 64463 56287
rect 32965 55913 32999 55947
rect 49249 55913 49283 55947
rect 64245 55913 64279 55947
rect 33793 55709 33827 55743
rect 48697 55709 48731 55743
rect 49157 55709 49191 55743
rect 63693 55709 63727 55743
rect 64337 55709 64371 55743
rect 64889 55709 64923 55743
rect 65625 55709 65659 55743
rect 63601 55573 63635 55607
rect 64981 55573 65015 55607
rect 50537 55301 50571 55335
rect 65165 55301 65199 55335
rect 66821 55301 66855 55335
rect 33517 55233 33551 55267
rect 35357 55233 35391 55267
rect 48697 55233 48731 55267
rect 64981 55233 65015 55267
rect 35173 55165 35207 55199
rect 48881 55165 48915 55199
rect 63693 55029 63727 55063
rect 33609 54825 33643 54859
rect 34805 54825 34839 54859
rect 48697 54825 48731 54859
rect 63233 54689 63267 54723
rect 63417 54689 63451 54723
rect 65073 54689 65107 54723
rect 33701 54621 33735 54655
rect 34897 54621 34931 54655
rect 48605 54621 48639 54655
rect 40785 52853 40819 52887
rect 40693 52513 40727 52547
rect 41153 52513 41187 52547
rect 40877 52377 40911 52411
rect 40877 52105 40911 52139
rect 40785 51969 40819 52003
rect 31585 51901 31619 51935
rect 32137 51901 32171 51935
rect 32321 51901 32355 51935
rect 32597 51901 32631 51935
rect 51089 51765 51123 51799
rect 31861 51561 31895 51595
rect 50997 51425 51031 51459
rect 52837 51425 52871 51459
rect 31769 51357 31803 51391
rect 51181 51289 51215 51323
rect 50813 51017 50847 51051
rect 50721 50881 50755 50915
rect 24501 50677 24535 50711
rect 24869 50337 24903 50371
rect 24409 50269 24443 50303
rect 24593 50201 24627 50235
rect 24869 49929 24903 49963
rect 24961 49793 24995 49827
rect 54217 49181 54251 49215
rect 53481 48705 53515 48739
rect 54125 48705 54159 48739
rect 53573 48637 53607 48671
rect 54309 48637 54343 48671
rect 55965 48637 55999 48671
rect 21005 48501 21039 48535
rect 22661 48161 22695 48195
rect 20821 48025 20855 48059
rect 22477 48025 22511 48059
rect 21925 47753 21959 47787
rect 49433 47685 49467 47719
rect 22017 47617 22051 47651
rect 47041 47549 47075 47583
rect 47593 47549 47627 47583
rect 47777 47549 47811 47583
rect 61945 47413 61979 47447
rect 46949 47209 46983 47243
rect 57897 47073 57931 47107
rect 59737 47073 59771 47107
rect 61945 47073 61979 47107
rect 63785 47073 63819 47107
rect 46857 47005 46891 47039
rect 57253 47005 57287 47039
rect 57345 46937 57379 46971
rect 58081 46937 58115 46971
rect 62129 46937 62163 46971
rect 61761 46665 61795 46699
rect 57989 46529 58023 46563
rect 61669 46529 61703 46563
rect 42441 46325 42475 46359
rect 41981 45985 42015 46019
rect 42441 45985 42475 46019
rect 41337 45917 41371 45951
rect 61025 45917 61059 45951
rect 41429 45849 41463 45883
rect 42165 45849 42199 45883
rect 62497 45509 62531 45543
rect 60657 45441 60691 45475
rect 60841 45373 60875 45407
rect 60657 45033 60691 45067
rect 60565 44829 60599 44863
rect 60473 43741 60507 43775
rect 60289 43265 60323 43299
rect 60473 43197 60507 43231
rect 62037 43197 62071 43231
rect 16865 43061 16899 43095
rect 34161 43061 34195 43095
rect 45109 43061 45143 43095
rect 52745 43061 52779 43095
rect 60565 42857 60599 42891
rect 35173 42721 35207 42755
rect 45017 42721 45051 42755
rect 46857 42721 46891 42755
rect 52193 42721 52227 42755
rect 16773 42653 16807 42687
rect 34713 42653 34747 42687
rect 51549 42653 51583 42687
rect 60473 42653 60507 42687
rect 16957 42585 16991 42619
rect 18613 42585 18647 42619
rect 34897 42585 34931 42619
rect 45201 42585 45235 42619
rect 51641 42585 51675 42619
rect 52377 42585 52411 42619
rect 54033 42585 54067 42619
rect 16957 42313 16991 42347
rect 34621 42313 34655 42347
rect 45017 42313 45051 42347
rect 16865 42177 16899 42211
rect 34713 42177 34747 42211
rect 44925 42177 44959 42211
rect 57897 41973 57931 42007
rect 57437 41633 57471 41667
rect 59093 41633 59127 41667
rect 56793 41565 56827 41599
rect 56885 41497 56919 41531
rect 57621 41497 57655 41531
rect 9873 39797 9907 39831
rect 9781 39457 9815 39491
rect 10241 39457 10275 39491
rect 33057 39389 33091 39423
rect 9965 39321 9999 39355
rect 10425 39049 10459 39083
rect 64797 38981 64831 39015
rect 65533 38981 65567 39015
rect 10517 38913 10551 38947
rect 32965 38913 32999 38947
rect 64705 38913 64739 38947
rect 33149 38845 33183 38879
rect 34805 38845 34839 38879
rect 65349 38845 65383 38879
rect 67189 38845 67223 38879
rect 32965 38505 32999 38539
rect 65625 38505 65659 38539
rect 32873 38301 32907 38335
rect 37381 37621 37415 37655
rect 61669 37621 61703 37655
rect 37381 37281 37415 37315
rect 61669 37281 61703 37315
rect 63509 37281 63543 37315
rect 35357 37213 35391 37247
rect 39221 37213 39255 37247
rect 61025 37213 61059 37247
rect 32413 37145 32447 37179
rect 37565 37145 37599 37179
rect 61117 37145 61151 37179
rect 61853 37145 61887 37179
rect 32505 37077 32539 37111
rect 35541 37077 35575 37111
rect 36645 36873 36679 36907
rect 35449 36805 35483 36839
rect 37933 36805 37967 36839
rect 38945 36805 38979 36839
rect 40325 36805 40359 36839
rect 33149 36737 33183 36771
rect 34069 36737 34103 36771
rect 35817 36737 35851 36771
rect 36553 36737 36587 36771
rect 37381 36737 37415 36771
rect 38577 36737 38611 36771
rect 39773 36737 39807 36771
rect 64797 36737 64831 36771
rect 13461 36669 13495 36703
rect 13921 36669 13955 36703
rect 14105 36669 14139 36703
rect 14381 36669 14415 36703
rect 34437 36669 34471 36703
rect 33425 36533 33459 36567
rect 64889 36533 64923 36567
rect 65625 36533 65659 36567
rect 14197 36329 14231 36363
rect 38117 36193 38151 36227
rect 65625 36193 65659 36227
rect 65809 36193 65843 36227
rect 6377 36125 6411 36159
rect 14289 36125 14323 36159
rect 32413 36125 32447 36159
rect 33517 36125 33551 36159
rect 33793 36125 33827 36159
rect 36093 36125 36127 36159
rect 36553 36125 36587 36159
rect 37565 36125 37599 36159
rect 45385 36125 45419 36159
rect 32965 36057 32999 36091
rect 35265 36057 35299 36091
rect 67465 36057 67499 36091
rect 36737 35989 36771 36023
rect 34529 35717 34563 35751
rect 47041 35717 47075 35751
rect 6377 35649 6411 35683
rect 32873 35649 32907 35683
rect 33977 35649 34011 35683
rect 35909 35649 35943 35683
rect 44557 35649 44591 35683
rect 45201 35649 45235 35683
rect 6561 35581 6595 35615
rect 6837 35581 6871 35615
rect 32597 35581 32631 35615
rect 35357 35581 35391 35615
rect 44649 35581 44683 35615
rect 45385 35581 45419 35615
rect 6469 35241 6503 35275
rect 6561 35037 6595 35071
rect 35909 34561 35943 34595
rect 37381 34561 37415 34595
rect 35265 34493 35299 34527
rect 37933 34493 37967 34527
rect 24869 34357 24903 34391
rect 24869 34017 24903 34051
rect 25329 34017 25363 34051
rect 35449 34017 35483 34051
rect 36737 34017 36771 34051
rect 35725 33949 35759 33983
rect 37013 33949 37047 33983
rect 49249 33949 49283 33983
rect 55873 33949 55907 33983
rect 25053 33881 25087 33915
rect 25237 33609 25271 33643
rect 25329 33473 25363 33507
rect 41705 33473 41739 33507
rect 49157 33473 49191 33507
rect 55505 33473 55539 33507
rect 42441 33405 42475 33439
rect 42625 33405 42659 33439
rect 44281 33405 44315 33439
rect 49341 33405 49375 33439
rect 50997 33405 51031 33439
rect 55689 33405 55723 33439
rect 57345 33405 57379 33439
rect 41797 33337 41831 33371
rect 42257 33065 42291 33099
rect 49157 33065 49191 33099
rect 56149 33065 56183 33099
rect 49065 32861 49099 32895
rect 56241 32861 56275 32895
rect 44005 32453 44039 32487
rect 44741 32453 44775 32487
rect 43913 32385 43947 32419
rect 44557 32317 44591 32351
rect 45017 32317 45051 32351
rect 45017 31977 45051 32011
rect 5457 31773 5491 31807
rect 6561 31297 6595 31331
rect 38301 31297 38335 31331
rect 38853 31229 38887 31263
rect 6469 31093 6503 31127
rect 5457 30753 5491 30787
rect 5641 30753 5675 30787
rect 5917 30753 5951 30787
rect 32873 30753 32907 30787
rect 7849 30685 7883 30719
rect 19533 30685 19567 30719
rect 28089 30685 28123 30719
rect 33425 30685 33459 30719
rect 59737 30685 59771 30719
rect 60473 30685 60507 30719
rect 59829 30617 59863 30651
rect 60657 30617 60691 30651
rect 62313 30617 62347 30651
rect 7757 30209 7791 30243
rect 19441 30209 19475 30243
rect 26157 30209 26191 30243
rect 27997 30209 28031 30243
rect 60197 30209 60231 30243
rect 7941 30141 7975 30175
rect 8401 30141 8435 30175
rect 19625 30141 19659 30175
rect 20085 30141 20119 30175
rect 28181 30141 28215 30175
rect 28457 30141 28491 30175
rect 25513 30005 25547 30039
rect 26065 30005 26099 30039
rect 27537 30005 27571 30039
rect 51181 30005 51215 30039
rect 8309 29801 8343 29835
rect 19993 29801 20027 29835
rect 28365 29801 28399 29835
rect 25513 29665 25547 29699
rect 25697 29665 25731 29699
rect 25973 29665 26007 29699
rect 8401 29597 8435 29631
rect 20085 29597 20119 29631
rect 28457 29597 28491 29631
rect 50905 29597 50939 29631
rect 51549 29597 51583 29631
rect 51733 29529 51767 29563
rect 53389 29529 53423 29563
rect 50997 29461 51031 29495
rect 51549 29189 51583 29223
rect 27537 29121 27571 29155
rect 37381 29121 37415 29155
rect 39129 29121 39163 29155
rect 51457 29121 51491 29155
rect 27721 29053 27755 29087
rect 27997 29053 28031 29087
rect 37841 29053 37875 29087
rect 38853 29053 38887 29087
rect 50997 28985 51031 29019
rect 28089 28713 28123 28747
rect 51089 28577 51123 28611
rect 51273 28577 51307 28611
rect 28181 28509 28215 28543
rect 33609 28509 33643 28543
rect 61209 28509 61243 28543
rect 33149 28441 33183 28475
rect 52929 28441 52963 28475
rect 60657 28033 60691 28067
rect 49893 27965 49927 27999
rect 50353 27965 50387 27999
rect 50537 27965 50571 27999
rect 52193 27965 52227 27999
rect 60841 27965 60875 27999
rect 62497 27965 62531 27999
rect 50537 27625 50571 27659
rect 61209 27625 61243 27659
rect 50445 27421 50479 27455
rect 61301 27421 61335 27455
rect 33793 26877 33827 26911
rect 33977 26877 34011 26911
rect 34897 26877 34931 26911
rect 56425 26741 56459 26775
rect 58265 26741 58299 26775
rect 33793 26537 33827 26571
rect 34805 26537 34839 26571
rect 55781 26401 55815 26435
rect 58081 26401 58115 26435
rect 26157 26333 26191 26367
rect 34897 26333 34931 26367
rect 59921 26333 59955 26367
rect 55965 26265 55999 26299
rect 57621 26265 57655 26299
rect 58265 26265 58299 26299
rect 56425 25993 56459 26027
rect 58265 25993 58299 26027
rect 27169 25857 27203 25891
rect 56517 25857 56551 25891
rect 58173 25857 58207 25891
rect 27077 25653 27111 25687
rect 27537 25313 27571 25347
rect 27721 25313 27755 25347
rect 32689 25313 32723 25347
rect 12357 25245 12391 25279
rect 28181 25245 28215 25279
rect 32229 25245 32263 25279
rect 25881 25177 25915 25211
rect 32137 25109 32171 25143
rect 32321 24837 32355 24871
rect 12357 24769 12391 24803
rect 23673 24769 23707 24803
rect 28181 24769 28215 24803
rect 32137 24769 32171 24803
rect 12541 24701 12575 24735
rect 13093 24701 13127 24735
rect 28365 24701 28399 24735
rect 28641 24701 28675 24735
rect 32597 24701 32631 24735
rect 23029 24565 23063 24599
rect 23581 24565 23615 24599
rect 13001 24361 13035 24395
rect 28549 24361 28583 24395
rect 13093 24157 13127 24191
rect 28641 24157 28675 24191
rect 23213 23749 23247 23783
rect 23029 23681 23063 23715
rect 24685 23613 24719 23647
rect 51733 22661 51767 22695
rect 52929 22661 52963 22695
rect 51641 22593 51675 22627
rect 52745 22525 52779 22559
rect 54585 22525 54619 22559
rect 6561 22389 6595 22423
rect 9321 22389 9355 22423
rect 11805 22389 11839 22423
rect 56425 22389 56459 22423
rect 61853 22389 61887 22423
rect 52193 22185 52227 22219
rect 7573 22049 7607 22083
rect 9321 22049 9355 22083
rect 9505 22049 9539 22083
rect 9781 22049 9815 22083
rect 11713 22049 11747 22083
rect 13093 22049 13127 22083
rect 26617 22049 26651 22083
rect 56333 22049 56367 22083
rect 57897 22049 57931 22083
rect 61761 22049 61795 22083
rect 25513 21981 25547 22015
rect 26157 21981 26191 22015
rect 5733 21913 5767 21947
rect 7389 21913 7423 21947
rect 11897 21913 11931 21947
rect 25605 21913 25639 21947
rect 26341 21913 26375 21947
rect 56517 21913 56551 21947
rect 61945 21913 61979 21947
rect 63601 21913 63635 21947
rect 6469 21641 6503 21675
rect 9689 21641 9723 21675
rect 12081 21641 12115 21675
rect 56333 21641 56367 21675
rect 61761 21641 61795 21675
rect 6561 21505 6595 21539
rect 9781 21505 9815 21539
rect 12173 21505 12207 21539
rect 56241 21505 56275 21539
rect 61669 21505 61703 21539
rect 26249 21437 26283 21471
rect 27353 20961 27387 20995
rect 8953 20893 8987 20927
rect 27169 20893 27203 20927
rect 62681 20893 62715 20927
rect 8677 20417 8711 20451
rect 62221 20417 62255 20451
rect 63049 20417 63083 20451
rect 64889 20417 64923 20451
rect 8861 20349 8895 20383
rect 9137 20349 9171 20383
rect 62313 20349 62347 20383
rect 63233 20349 63267 20383
rect 9045 20009 9079 20043
rect 9137 19805 9171 19839
rect 27905 19329 27939 19363
rect 35173 19329 35207 19363
rect 35265 19193 35299 19227
rect 27997 19125 28031 19159
rect 28733 19125 28767 19159
rect 35817 19125 35851 19159
rect 28825 18785 28859 18819
rect 29009 18785 29043 18819
rect 35541 18785 35575 18819
rect 35725 18785 35759 18819
rect 37197 18785 37231 18819
rect 23857 18717 23891 18751
rect 24777 18717 24811 18751
rect 27169 18649 27203 18683
rect 24685 18581 24719 18615
rect 24317 18309 24351 18343
rect 24133 18241 24167 18275
rect 24593 18173 24627 18207
rect 38485 17697 38519 17731
rect 14105 17629 14139 17663
rect 36185 17629 36219 17663
rect 36829 17629 36863 17663
rect 58817 17629 58851 17663
rect 59461 17629 59495 17663
rect 36277 17561 36311 17595
rect 37013 17561 37047 17595
rect 58909 17493 58943 17527
rect 59369 17221 59403 17255
rect 13737 17153 13771 17187
rect 37289 17153 37323 17187
rect 59185 17153 59219 17187
rect 13921 17085 13955 17119
rect 14473 17085 14507 17119
rect 61025 17085 61059 17119
rect 14197 16745 14231 16779
rect 14289 16551 14323 16585
rect 23213 15453 23247 15487
rect 23857 15453 23891 15487
rect 62037 15453 62071 15487
rect 62865 15453 62899 15487
rect 23765 15317 23799 15351
rect 62129 15317 62163 15351
rect 23305 15045 23339 15079
rect 63233 15045 63267 15079
rect 23121 14977 23155 15011
rect 63049 14977 63083 15011
rect 23581 14909 23615 14943
rect 64797 14909 64831 14943
rect 15025 14365 15059 14399
rect 35725 14365 35759 14399
rect 36369 14365 36403 14399
rect 15117 14229 15151 14263
rect 35817 14229 35851 14263
rect 30665 13957 30699 13991
rect 30757 13889 30791 13923
rect 10701 13821 10735 13855
rect 31401 13821 31435 13855
rect 15025 13685 15059 13719
rect 10425 13345 10459 13379
rect 12265 13345 12299 13379
rect 14933 13345 14967 13379
rect 15117 13345 15151 13379
rect 15485 13345 15519 13379
rect 31953 13345 31987 13379
rect 32137 13345 32171 13379
rect 35633 13345 35667 13379
rect 35817 13345 35851 13379
rect 36093 13345 36127 13379
rect 12081 13209 12115 13243
rect 30297 13209 30331 13243
rect 11621 12937 11655 12971
rect 11713 12801 11747 12835
rect 9045 12597 9079 12631
rect 8309 12189 8343 12223
rect 9689 12189 9723 12223
rect 40233 12189 40267 12223
rect 41521 12189 41555 12223
rect 9597 12053 9631 12087
rect 41613 12053 41647 12087
rect 9229 11781 9263 11815
rect 8401 11713 8435 11747
rect 9045 11713 9079 11747
rect 40049 11713 40083 11747
rect 9781 11645 9815 11679
rect 40233 11645 40267 11679
rect 41889 11645 41923 11679
rect 8493 11509 8527 11543
rect 24409 11509 24443 11543
rect 42441 11509 42475 11543
rect 40141 11305 40175 11339
rect 8953 11169 8987 11203
rect 9137 11169 9171 11203
rect 9873 11169 9907 11203
rect 24409 11169 24443 11203
rect 24869 11169 24903 11203
rect 41705 11169 41739 11203
rect 41889 11169 41923 11203
rect 27537 11101 27571 11135
rect 40049 11101 40083 11135
rect 24593 11033 24627 11067
rect 43545 11033 43579 11067
rect 24777 10761 24811 10795
rect 10241 10625 10275 10659
rect 24869 10625 24903 10659
rect 27537 10625 27571 10659
rect 38209 10625 38243 10659
rect 44005 10625 44039 10659
rect 27721 10557 27755 10591
rect 29377 10557 29411 10591
rect 9597 10421 9631 10455
rect 10149 10421 10183 10455
rect 38301 10421 38335 10455
rect 38853 10421 38887 10455
rect 44097 10421 44131 10455
rect 44833 10421 44867 10455
rect 27905 10217 27939 10251
rect 9781 10081 9815 10115
rect 9965 10081 9999 10115
rect 10333 10081 10367 10115
rect 45017 10081 45051 10115
rect 45201 10081 45235 10115
rect 27997 10013 28031 10047
rect 46857 9945 46891 9979
rect 38301 9605 38335 9639
rect 38117 9469 38151 9503
rect 38669 9469 38703 9503
rect 47869 8245 47903 8279
rect 47777 7905 47811 7939
rect 47133 7837 47167 7871
rect 47225 7769 47259 7803
rect 47961 7769 47995 7803
rect 49617 7769 49651 7803
rect 10885 6749 10919 6783
rect 11345 6749 11379 6783
rect 11989 6749 12023 6783
rect 11437 6613 11471 6647
rect 11713 6341 11747 6375
rect 10793 6273 10827 6307
rect 11529 6273 11563 6307
rect 43361 6273 43395 6307
rect 12449 6205 12483 6239
rect 10885 6069 10919 6103
rect 43453 6069 43487 6103
rect 11161 5729 11195 5763
rect 11345 5729 11379 5763
rect 11621 5729 11655 5763
rect 43545 5661 43579 5695
rect 43637 5253 43671 5287
rect 43453 5185 43487 5219
rect 45293 5117 45327 5151
rect 12449 4981 12483 5015
rect 29561 4709 29595 4743
rect 13553 4641 13587 4675
rect 29009 4573 29043 4607
rect 11713 4505 11747 4539
rect 13369 4505 13403 4539
rect 12541 4233 12575 4267
rect 12449 4097 12483 4131
rect 28365 4097 28399 4131
rect 29009 4097 29043 4131
rect 29193 4029 29227 4063
rect 29653 4029 29687 4063
rect 28457 3961 28491 3995
rect 29561 3553 29595 3587
rect 28825 3485 28859 3519
rect 28917 3417 28951 3451
rect 29745 3417 29779 3451
rect 31401 3417 31435 3451
<< metal1 >>
rect 1104 69658 68816 69680
rect 1104 69606 19574 69658
rect 19626 69606 19638 69658
rect 19690 69606 19702 69658
rect 19754 69606 19766 69658
rect 19818 69606 19830 69658
rect 19882 69606 50294 69658
rect 50346 69606 50358 69658
rect 50410 69606 50422 69658
rect 50474 69606 50486 69658
rect 50538 69606 50550 69658
rect 50602 69606 68816 69658
rect 1104 69584 68816 69606
rect 62758 69164 62764 69216
rect 62816 69204 62822 69216
rect 66070 69204 66076 69216
rect 62816 69176 66076 69204
rect 62816 69164 62822 69176
rect 66070 69164 66076 69176
rect 66128 69164 66134 69216
rect 1104 69114 68816 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 34934 69114
rect 34986 69062 34998 69114
rect 35050 69062 35062 69114
rect 35114 69062 35126 69114
rect 35178 69062 35190 69114
rect 35242 69062 65654 69114
rect 65706 69062 65718 69114
rect 65770 69062 65782 69114
rect 65834 69062 65846 69114
rect 65898 69062 65910 69114
rect 65962 69062 68816 69114
rect 1104 69040 68816 69062
rect 52822 68960 52828 69012
rect 52880 69000 52886 69012
rect 56686 69000 56692 69012
rect 52880 68972 56692 69000
rect 52880 68960 52886 68972
rect 56686 68960 56692 68972
rect 56744 68960 56750 69012
rect 62022 68756 62028 68808
rect 62080 68796 62086 68808
rect 65334 68796 65340 68808
rect 62080 68768 65340 68796
rect 62080 68756 62086 68768
rect 65334 68756 65340 68768
rect 65392 68756 65398 68808
rect 1104 68570 68816 68592
rect 1104 68518 19574 68570
rect 19626 68518 19638 68570
rect 19690 68518 19702 68570
rect 19754 68518 19766 68570
rect 19818 68518 19830 68570
rect 19882 68518 50294 68570
rect 50346 68518 50358 68570
rect 50410 68518 50422 68570
rect 50474 68518 50486 68570
rect 50538 68518 50550 68570
rect 50602 68518 68816 68570
rect 1104 68496 68816 68518
rect 1946 68280 1952 68332
rect 2004 68320 2010 68332
rect 15838 68320 15844 68332
rect 2004 68292 15844 68320
rect 2004 68280 2010 68292
rect 15838 68280 15844 68292
rect 15896 68280 15902 68332
rect 21266 68280 21272 68332
rect 21324 68320 21330 68332
rect 35342 68320 35348 68332
rect 21324 68292 35348 68320
rect 21324 68280 21330 68292
rect 35342 68280 35348 68292
rect 35400 68280 35406 68332
rect 50614 68280 50620 68332
rect 50672 68320 50678 68332
rect 66990 68320 66996 68332
rect 50672 68292 66996 68320
rect 50672 68280 50678 68292
rect 66990 68280 66996 68292
rect 67048 68280 67054 68332
rect 49418 68144 49424 68196
rect 49476 68184 49482 68196
rect 54110 68184 54116 68196
rect 49476 68156 54116 68184
rect 49476 68144 49482 68156
rect 54110 68144 54116 68156
rect 54168 68144 54174 68196
rect 46842 68076 46848 68128
rect 46900 68116 46906 68128
rect 51534 68116 51540 68128
rect 46900 68088 51540 68116
rect 46900 68076 46906 68088
rect 51534 68076 51540 68088
rect 51592 68076 51598 68128
rect 1104 68026 68816 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 34934 68026
rect 34986 67974 34998 68026
rect 35050 67974 35062 68026
rect 35114 67974 35126 68026
rect 35178 67974 35190 68026
rect 35242 67974 65654 68026
rect 65706 67974 65718 68026
rect 65770 67974 65782 68026
rect 65834 67974 65846 68026
rect 65898 67974 65910 68026
rect 65962 67974 68816 68026
rect 1104 67952 68816 67974
rect 48958 67872 48964 67924
rect 49016 67912 49022 67924
rect 49878 67912 49884 67924
rect 49016 67884 49884 67912
rect 49016 67872 49022 67884
rect 49878 67872 49884 67884
rect 49936 67872 49942 67924
rect 19978 67736 19984 67788
rect 20036 67776 20042 67788
rect 21266 67776 21272 67788
rect 20036 67748 21272 67776
rect 20036 67736 20042 67748
rect 21266 67736 21272 67748
rect 21324 67736 21330 67788
rect 1104 67482 68816 67504
rect 1104 67430 19574 67482
rect 19626 67430 19638 67482
rect 19690 67430 19702 67482
rect 19754 67430 19766 67482
rect 19818 67430 19830 67482
rect 19882 67430 50294 67482
rect 50346 67430 50358 67482
rect 50410 67430 50422 67482
rect 50474 67430 50486 67482
rect 50538 67430 50550 67482
rect 50602 67430 68816 67482
rect 1104 67408 68816 67430
rect 1104 66938 68816 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 68816 66938
rect 1104 66864 68816 66886
rect 1104 66394 68816 66416
rect 1104 66342 19574 66394
rect 19626 66342 19638 66394
rect 19690 66342 19702 66394
rect 19754 66342 19766 66394
rect 19818 66342 19830 66394
rect 19882 66342 50294 66394
rect 50346 66342 50358 66394
rect 50410 66342 50422 66394
rect 50474 66342 50486 66394
rect 50538 66342 50550 66394
rect 50602 66342 68816 66394
rect 1104 66320 68816 66342
rect 39206 66240 39212 66292
rect 39264 66280 39270 66292
rect 65334 66280 65340 66292
rect 39264 66252 65340 66280
rect 39264 66240 39270 66252
rect 65334 66240 65340 66252
rect 65392 66240 65398 66292
rect 1394 66144 1400 66156
rect 1355 66116 1400 66144
rect 1394 66104 1400 66116
rect 1452 66104 1458 66156
rect 1578 66076 1584 66088
rect 1539 66048 1584 66076
rect 1578 66036 1584 66048
rect 1636 66036 1642 66088
rect 1104 65850 68816 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 68816 65850
rect 1104 65776 68816 65798
rect 1104 65306 68816 65328
rect 1104 65254 19574 65306
rect 19626 65254 19638 65306
rect 19690 65254 19702 65306
rect 19754 65254 19766 65306
rect 19818 65254 19830 65306
rect 19882 65254 50294 65306
rect 50346 65254 50358 65306
rect 50410 65254 50422 65306
rect 50474 65254 50486 65306
rect 50538 65254 50550 65306
rect 50602 65254 68816 65306
rect 1104 65232 68816 65254
rect 1104 64762 68816 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 34934 64762
rect 34986 64710 34998 64762
rect 35050 64710 35062 64762
rect 35114 64710 35126 64762
rect 35178 64710 35190 64762
rect 35242 64710 65654 64762
rect 65706 64710 65718 64762
rect 65770 64710 65782 64762
rect 65834 64710 65846 64762
rect 65898 64710 65910 64762
rect 65962 64710 68816 64762
rect 1104 64688 68816 64710
rect 19426 64404 19432 64456
rect 19484 64444 19490 64456
rect 19797 64447 19855 64453
rect 19797 64444 19809 64447
rect 19484 64416 19809 64444
rect 19484 64404 19490 64416
rect 19797 64413 19809 64416
rect 19843 64413 19855 64447
rect 19797 64407 19855 64413
rect 1104 64218 68816 64240
rect 1104 64166 19574 64218
rect 19626 64166 19638 64218
rect 19690 64166 19702 64218
rect 19754 64166 19766 64218
rect 19818 64166 19830 64218
rect 19882 64166 50294 64218
rect 50346 64166 50358 64218
rect 50410 64166 50422 64218
rect 50474 64166 50486 64218
rect 50538 64166 50550 64218
rect 50602 64166 68816 64218
rect 1104 64144 68816 64166
rect 21266 64036 21272 64048
rect 21227 64008 21272 64036
rect 21266 63996 21272 64008
rect 21324 63996 21330 64048
rect 19426 63968 19432 63980
rect 19387 63940 19432 63968
rect 19426 63928 19432 63940
rect 19484 63928 19490 63980
rect 19613 63903 19671 63909
rect 19613 63869 19625 63903
rect 19659 63900 19671 63903
rect 20162 63900 20168 63912
rect 19659 63872 20168 63900
rect 19659 63869 19671 63872
rect 19613 63863 19671 63869
rect 20162 63860 20168 63872
rect 20220 63860 20226 63912
rect 18969 63767 19027 63773
rect 18969 63733 18981 63767
rect 19015 63764 19027 63767
rect 19334 63764 19340 63776
rect 19015 63736 19340 63764
rect 19015 63733 19027 63736
rect 18969 63727 19027 63733
rect 19334 63724 19340 63736
rect 19392 63724 19398 63776
rect 1104 63674 68816 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 34934 63674
rect 34986 63622 34998 63674
rect 35050 63622 35062 63674
rect 35114 63622 35126 63674
rect 35178 63622 35190 63674
rect 35242 63622 65654 63674
rect 65706 63622 65718 63674
rect 65770 63622 65782 63674
rect 65834 63622 65846 63674
rect 65898 63622 65910 63674
rect 65962 63622 68816 63674
rect 1104 63600 68816 63622
rect 15838 63452 15844 63504
rect 15896 63492 15902 63504
rect 15896 63464 19840 63492
rect 15896 63452 15902 63464
rect 19334 63424 19340 63436
rect 19295 63396 19340 63424
rect 19334 63384 19340 63396
rect 19392 63384 19398 63436
rect 19812 63433 19840 63464
rect 19797 63427 19855 63433
rect 19797 63393 19809 63427
rect 19843 63393 19855 63427
rect 19797 63387 19855 63393
rect 43346 63356 43352 63368
rect 43307 63328 43352 63356
rect 43346 63316 43352 63328
rect 43404 63316 43410 63368
rect 43622 63316 43628 63368
rect 43680 63356 43686 63368
rect 43993 63359 44051 63365
rect 43993 63356 44005 63359
rect 43680 63328 44005 63356
rect 43680 63316 43686 63328
rect 43993 63325 44005 63328
rect 44039 63325 44051 63359
rect 43993 63319 44051 63325
rect 19521 63291 19579 63297
rect 19521 63257 19533 63291
rect 19567 63257 19579 63291
rect 19521 63251 19579 63257
rect 19426 63180 19432 63232
rect 19484 63220 19490 63232
rect 19536 63220 19564 63251
rect 19484 63192 19564 63220
rect 43441 63223 43499 63229
rect 19484 63180 19490 63192
rect 43441 63189 43453 63223
rect 43487 63220 43499 63223
rect 43806 63220 43812 63232
rect 43487 63192 43812 63220
rect 43487 63189 43499 63192
rect 43441 63183 43499 63189
rect 43806 63180 43812 63192
rect 43864 63180 43870 63232
rect 1104 63130 68816 63152
rect 1104 63078 19574 63130
rect 19626 63078 19638 63130
rect 19690 63078 19702 63130
rect 19754 63078 19766 63130
rect 19818 63078 19830 63130
rect 19882 63078 50294 63130
rect 50346 63078 50358 63130
rect 50410 63078 50422 63130
rect 50474 63078 50486 63130
rect 50538 63078 50550 63130
rect 50602 63078 68816 63130
rect 1104 63056 68816 63078
rect 19426 62976 19432 63028
rect 19484 63016 19490 63028
rect 19521 63019 19579 63025
rect 19521 63016 19533 63019
rect 19484 62988 19533 63016
rect 19484 62976 19490 62988
rect 19521 62985 19533 62988
rect 19567 62985 19579 63019
rect 20162 63016 20168 63028
rect 20123 62988 20168 63016
rect 19521 62979 19579 62985
rect 20162 62976 20168 62988
rect 20220 62976 20226 63028
rect 43806 62948 43812 62960
rect 43767 62920 43812 62948
rect 43806 62908 43812 62920
rect 43864 62908 43870 62960
rect 19613 62883 19671 62889
rect 19613 62849 19625 62883
rect 19659 62880 19671 62883
rect 20257 62883 20315 62889
rect 20257 62880 20269 62883
rect 19659 62852 20269 62880
rect 19659 62849 19671 62852
rect 19613 62843 19671 62849
rect 20257 62849 20269 62852
rect 20303 62880 20315 62883
rect 43346 62880 43352 62892
rect 20303 62852 43352 62880
rect 20303 62849 20315 62852
rect 20257 62843 20315 62849
rect 43346 62840 43352 62852
rect 43404 62840 43410 62892
rect 43622 62880 43628 62892
rect 43583 62852 43628 62880
rect 43622 62840 43628 62852
rect 43680 62840 43686 62892
rect 45465 62815 45523 62821
rect 45465 62781 45477 62815
rect 45511 62812 45523 62815
rect 48958 62812 48964 62824
rect 45511 62784 48964 62812
rect 45511 62781 45523 62784
rect 45465 62775 45523 62781
rect 48958 62772 48964 62784
rect 49016 62772 49022 62824
rect 1104 62586 68816 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 34934 62586
rect 34986 62534 34998 62586
rect 35050 62534 35062 62586
rect 35114 62534 35126 62586
rect 35178 62534 35190 62586
rect 35242 62534 65654 62586
rect 65706 62534 65718 62586
rect 65770 62534 65782 62586
rect 65834 62534 65846 62586
rect 65898 62534 65910 62586
rect 65962 62534 68816 62586
rect 1104 62512 68816 62534
rect 32766 62228 32772 62280
rect 32824 62268 32830 62280
rect 37093 62271 37151 62277
rect 32824 62240 32869 62268
rect 32824 62228 32830 62240
rect 37093 62237 37105 62271
rect 37139 62268 37151 62271
rect 37274 62268 37280 62280
rect 37139 62240 37280 62268
rect 37139 62237 37151 62240
rect 37093 62231 37151 62237
rect 37274 62228 37280 62240
rect 37332 62228 37338 62280
rect 5534 62160 5540 62212
rect 5592 62200 5598 62212
rect 30929 62203 30987 62209
rect 30929 62200 30941 62203
rect 5592 62172 30941 62200
rect 5592 62160 5598 62172
rect 30929 62169 30941 62172
rect 30975 62169 30987 62203
rect 32582 62200 32588 62212
rect 32543 62172 32588 62200
rect 30929 62163 30987 62169
rect 32582 62160 32588 62172
rect 32640 62160 32646 62212
rect 1104 62042 68816 62064
rect 1104 61990 19574 62042
rect 19626 61990 19638 62042
rect 19690 61990 19702 62042
rect 19754 61990 19766 62042
rect 19818 61990 19830 62042
rect 19882 61990 50294 62042
rect 50346 61990 50358 62042
rect 50410 61990 50422 62042
rect 50474 61990 50486 62042
rect 50538 61990 50550 62042
rect 50602 61990 68816 62042
rect 1104 61968 68816 61990
rect 32217 61931 32275 61937
rect 32217 61897 32229 61931
rect 32263 61928 32275 61931
rect 32582 61928 32588 61940
rect 32263 61900 32588 61928
rect 32263 61897 32275 61900
rect 32217 61891 32275 61897
rect 32582 61888 32588 61900
rect 32640 61888 32646 61940
rect 54110 61860 54116 61872
rect 36556 61832 54116 61860
rect 32309 61795 32367 61801
rect 32309 61761 32321 61795
rect 32355 61792 32367 61795
rect 35618 61792 35624 61804
rect 32355 61764 35624 61792
rect 32355 61761 32367 61764
rect 32309 61755 32367 61761
rect 35618 61752 35624 61764
rect 35676 61792 35682 61804
rect 36556 61801 36584 61832
rect 54110 61820 54116 61832
rect 54168 61820 54174 61872
rect 36541 61795 36599 61801
rect 36541 61792 36553 61795
rect 35676 61764 36553 61792
rect 35676 61752 35682 61764
rect 36541 61761 36553 61764
rect 36587 61761 36599 61795
rect 37274 61792 37280 61804
rect 37235 61764 37280 61792
rect 36541 61755 36599 61761
rect 37274 61752 37280 61764
rect 37332 61752 37338 61804
rect 31205 61727 31263 61733
rect 31205 61693 31217 61727
rect 31251 61724 31263 61727
rect 32766 61724 32772 61736
rect 31251 61696 32772 61724
rect 31251 61693 31263 61696
rect 31205 61687 31263 61693
rect 32766 61684 32772 61696
rect 32824 61684 32830 61736
rect 36633 61727 36691 61733
rect 36633 61693 36645 61727
rect 36679 61724 36691 61727
rect 37461 61727 37519 61733
rect 37461 61724 37473 61727
rect 36679 61696 37473 61724
rect 36679 61693 36691 61696
rect 36633 61687 36691 61693
rect 37461 61693 37473 61696
rect 37507 61693 37519 61727
rect 37461 61687 37519 61693
rect 37737 61727 37795 61733
rect 37737 61693 37749 61727
rect 37783 61693 37795 61727
rect 37737 61687 37795 61693
rect 37366 61616 37372 61668
rect 37424 61656 37430 61668
rect 37752 61656 37780 61687
rect 37424 61628 37780 61656
rect 37424 61616 37430 61628
rect 45830 61548 45836 61600
rect 45888 61588 45894 61600
rect 45925 61591 45983 61597
rect 45925 61588 45937 61591
rect 45888 61560 45937 61588
rect 45888 61548 45894 61560
rect 45925 61557 45937 61560
rect 45971 61557 45983 61591
rect 45925 61551 45983 61557
rect 54757 61591 54815 61597
rect 54757 61557 54769 61591
rect 54803 61588 54815 61591
rect 55306 61588 55312 61600
rect 54803 61560 55312 61588
rect 54803 61557 54815 61560
rect 54757 61551 54815 61557
rect 55306 61548 55312 61560
rect 55364 61548 55370 61600
rect 1104 61498 68816 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 65654 61498
rect 65706 61446 65718 61498
rect 65770 61446 65782 61498
rect 65834 61446 65846 61498
rect 65898 61446 65910 61498
rect 65962 61446 68816 61498
rect 1104 61424 68816 61446
rect 45554 61276 45560 61328
rect 45612 61316 45618 61328
rect 45612 61288 46336 61316
rect 45612 61276 45618 61288
rect 45830 61248 45836 61260
rect 45791 61220 45836 61248
rect 45830 61208 45836 61220
rect 45888 61208 45894 61260
rect 46308 61257 46336 61288
rect 46293 61251 46351 61257
rect 46293 61217 46305 61251
rect 46339 61217 46351 61251
rect 55306 61248 55312 61260
rect 55267 61220 55312 61248
rect 46293 61211 46351 61217
rect 55306 61208 55312 61220
rect 55364 61208 55370 61260
rect 54110 61180 54116 61192
rect 54071 61152 54116 61180
rect 54110 61140 54116 61152
rect 54168 61140 54174 61192
rect 46014 61112 46020 61124
rect 45975 61084 46020 61112
rect 46014 61072 46020 61084
rect 46072 61072 46078 61124
rect 54205 61115 54263 61121
rect 54205 61081 54217 61115
rect 54251 61112 54263 61115
rect 55493 61115 55551 61121
rect 55493 61112 55505 61115
rect 54251 61084 55505 61112
rect 54251 61081 54263 61084
rect 54205 61075 54263 61081
rect 55493 61081 55505 61084
rect 55539 61081 55551 61115
rect 55493 61075 55551 61081
rect 57149 61115 57207 61121
rect 57149 61081 57161 61115
rect 57195 61112 57207 61115
rect 64874 61112 64880 61124
rect 57195 61084 64880 61112
rect 57195 61081 57207 61084
rect 57149 61075 57207 61081
rect 64874 61072 64880 61084
rect 64932 61072 64938 61124
rect 1104 60954 68816 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 68816 60954
rect 1104 60880 68816 60902
rect 46014 60840 46020 60852
rect 45975 60812 46020 60840
rect 46014 60800 46020 60812
rect 46072 60800 46078 60852
rect 3418 60732 3424 60784
rect 3476 60772 3482 60784
rect 24854 60772 24860 60784
rect 3476 60744 24860 60772
rect 3476 60732 3482 60744
rect 24854 60732 24860 60744
rect 24912 60732 24918 60784
rect 45922 60704 45928 60716
rect 45883 60676 45928 60704
rect 45922 60664 45928 60676
rect 45980 60664 45986 60716
rect 1104 60410 68816 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 65654 60410
rect 65706 60358 65718 60410
rect 65770 60358 65782 60410
rect 65834 60358 65846 60410
rect 65898 60358 65910 60410
rect 65962 60358 68816 60410
rect 1104 60336 68816 60358
rect 26513 60095 26571 60101
rect 26513 60061 26525 60095
rect 26559 60092 26571 60095
rect 26970 60092 26976 60104
rect 26559 60064 26976 60092
rect 26559 60061 26571 60064
rect 26513 60055 26571 60061
rect 26970 60052 26976 60064
rect 27028 60052 27034 60104
rect 35526 60052 35532 60104
rect 35584 60092 35590 60104
rect 35621 60095 35679 60101
rect 35621 60092 35633 60095
rect 35584 60064 35633 60092
rect 35584 60052 35590 60064
rect 35621 60061 35633 60064
rect 35667 60061 35679 60095
rect 35621 60055 35679 60061
rect 54846 60052 54852 60104
rect 54904 60092 54910 60104
rect 55309 60095 55367 60101
rect 55309 60092 55321 60095
rect 54904 60064 55321 60092
rect 54904 60052 54910 60064
rect 55309 60061 55321 60064
rect 55355 60061 55367 60095
rect 55309 60055 55367 60061
rect 1104 59866 68816 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 68816 59866
rect 1104 59792 68816 59814
rect 54297 59687 54355 59693
rect 26252 59656 35894 59684
rect 26252 59628 26280 59656
rect 26234 59576 26240 59628
rect 26292 59616 26298 59628
rect 26970 59616 26976 59628
rect 26292 59588 26385 59616
rect 26931 59588 26976 59616
rect 26292 59576 26298 59588
rect 26970 59576 26976 59588
rect 27028 59576 27034 59628
rect 26329 59551 26387 59557
rect 26329 59517 26341 59551
rect 26375 59548 26387 59551
rect 27157 59551 27215 59557
rect 27157 59548 27169 59551
rect 26375 59520 27169 59548
rect 26375 59517 26387 59520
rect 26329 59511 26387 59517
rect 27157 59517 27169 59520
rect 27203 59517 27215 59551
rect 27157 59511 27215 59517
rect 27433 59551 27491 59557
rect 27433 59517 27445 59551
rect 27479 59517 27491 59551
rect 27433 59511 27491 59517
rect 24854 59440 24860 59492
rect 24912 59480 24918 59492
rect 27448 59480 27476 59511
rect 24912 59452 27476 59480
rect 35866 59480 35894 59656
rect 54297 59653 54309 59687
rect 54343 59684 54355 59687
rect 55033 59687 55091 59693
rect 55033 59684 55045 59687
rect 54343 59656 55045 59684
rect 54343 59653 54355 59656
rect 54297 59647 54355 59653
rect 55033 59653 55045 59656
rect 55079 59653 55091 59687
rect 55033 59647 55091 59653
rect 56689 59687 56747 59693
rect 56689 59653 56701 59687
rect 56735 59684 56747 59687
rect 62758 59684 62764 59696
rect 56735 59656 62764 59684
rect 56735 59653 56747 59656
rect 56689 59647 56747 59653
rect 62758 59644 62764 59656
rect 62816 59644 62822 59696
rect 45922 59616 45928 59628
rect 45526 59588 45928 59616
rect 45526 59480 45554 59588
rect 45922 59576 45928 59588
rect 45980 59616 45986 59628
rect 54205 59619 54263 59625
rect 54205 59616 54217 59619
rect 45980 59588 54217 59616
rect 45980 59576 45986 59588
rect 54205 59585 54217 59588
rect 54251 59585 54263 59619
rect 54846 59616 54852 59628
rect 54807 59588 54852 59616
rect 54205 59579 54263 59585
rect 54846 59576 54852 59588
rect 54904 59576 54910 59628
rect 35866 59452 45554 59480
rect 24912 59440 24918 59452
rect 1104 59322 68816 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 65654 59322
rect 65706 59270 65718 59322
rect 65770 59270 65782 59322
rect 65834 59270 65846 59322
rect 65898 59270 65910 59322
rect 65962 59270 68816 59322
rect 1104 59248 68816 59270
rect 35526 59072 35532 59084
rect 35487 59044 35532 59072
rect 35526 59032 35532 59044
rect 35584 59032 35590 59084
rect 37182 59072 37188 59084
rect 37143 59044 37188 59072
rect 37182 59032 37188 59044
rect 37240 59032 37246 59084
rect 35710 58936 35716 58948
rect 35671 58908 35716 58936
rect 35710 58896 35716 58908
rect 35768 58896 35774 58948
rect 1104 58778 68816 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 68816 58778
rect 1104 58704 68816 58726
rect 35710 58664 35716 58676
rect 35671 58636 35716 58664
rect 35710 58624 35716 58636
rect 35768 58624 35774 58676
rect 66070 58556 66076 58608
rect 66128 58596 66134 58608
rect 66165 58599 66223 58605
rect 66165 58596 66177 58599
rect 66128 58568 66177 58596
rect 66128 58556 66134 58568
rect 66165 58565 66177 58568
rect 66211 58565 66223 58599
rect 66165 58559 66223 58565
rect 35434 58488 35440 58540
rect 35492 58528 35498 58540
rect 35621 58531 35679 58537
rect 35621 58528 35633 58531
rect 35492 58500 35633 58528
rect 35492 58488 35498 58500
rect 35621 58497 35633 58500
rect 35667 58497 35679 58531
rect 35621 58491 35679 58497
rect 37461 58531 37519 58537
rect 37461 58497 37473 58531
rect 37507 58528 37519 58531
rect 40310 58528 40316 58540
rect 37507 58500 40316 58528
rect 37507 58497 37519 58500
rect 37461 58491 37519 58497
rect 40310 58488 40316 58500
rect 40368 58488 40374 58540
rect 64325 58463 64383 58469
rect 64325 58429 64337 58463
rect 64371 58429 64383 58463
rect 64506 58460 64512 58472
rect 64467 58432 64512 58460
rect 64325 58423 64383 58429
rect 36541 58395 36599 58401
rect 36541 58361 36553 58395
rect 36587 58392 36599 58395
rect 38102 58392 38108 58404
rect 36587 58364 38108 58392
rect 36587 58361 36599 58364
rect 36541 58355 36599 58361
rect 38102 58352 38108 58364
rect 38160 58352 38166 58404
rect 64340 58392 64368 58423
rect 64506 58420 64512 58432
rect 64564 58420 64570 58472
rect 65518 58392 65524 58404
rect 64340 58364 65524 58392
rect 65518 58352 65524 58364
rect 65576 58352 65582 58404
rect 37369 58327 37427 58333
rect 37369 58293 37381 58327
rect 37415 58324 37427 58327
rect 37918 58324 37924 58336
rect 37415 58296 37924 58324
rect 37415 58293 37427 58296
rect 37369 58287 37427 58293
rect 37918 58284 37924 58296
rect 37976 58284 37982 58336
rect 1104 58234 68816 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 65654 58234
rect 65706 58182 65718 58234
rect 65770 58182 65782 58234
rect 65834 58182 65846 58234
rect 65898 58182 65910 58234
rect 65962 58182 68816 58234
rect 1104 58160 68816 58182
rect 64506 58080 64512 58132
rect 64564 58120 64570 58132
rect 64693 58123 64751 58129
rect 64693 58120 64705 58123
rect 64564 58092 64705 58120
rect 64564 58080 64570 58092
rect 64693 58089 64705 58092
rect 64739 58089 64751 58123
rect 64693 58083 64751 58089
rect 65518 58080 65524 58132
rect 65576 58120 65582 58132
rect 65613 58123 65671 58129
rect 65613 58120 65625 58123
rect 65576 58092 65625 58120
rect 65576 58080 65582 58092
rect 65613 58089 65625 58092
rect 65659 58089 65671 58123
rect 65613 58083 65671 58089
rect 37918 57984 37924 57996
rect 37879 57956 37924 57984
rect 37918 57944 37924 57956
rect 37976 57944 37982 57996
rect 40310 57944 40316 57996
rect 40368 57984 40374 57996
rect 63678 57984 63684 57996
rect 40368 57956 63684 57984
rect 40368 57944 40374 57956
rect 63678 57944 63684 57956
rect 63736 57984 63742 57996
rect 63736 57956 64000 57984
rect 63736 57944 63742 57956
rect 34698 57916 34704 57928
rect 34659 57888 34704 57916
rect 34698 57876 34704 57888
rect 34756 57876 34762 57928
rect 35342 57876 35348 57928
rect 35400 57916 35406 57928
rect 36265 57919 36323 57925
rect 36265 57916 36277 57919
rect 35400 57888 36277 57916
rect 35400 57876 35406 57888
rect 36265 57885 36277 57888
rect 36311 57885 36323 57919
rect 36265 57879 36323 57885
rect 38102 57876 38108 57928
rect 38160 57916 38166 57928
rect 63494 57916 63500 57928
rect 38160 57888 38205 57916
rect 63455 57888 63500 57916
rect 38160 57876 38166 57888
rect 63494 57876 63500 57888
rect 63552 57876 63558 57928
rect 63972 57925 64000 57956
rect 63957 57919 64015 57925
rect 63957 57885 63969 57919
rect 64003 57916 64015 57919
rect 64601 57919 64659 57925
rect 64601 57916 64613 57919
rect 64003 57888 64613 57916
rect 64003 57885 64015 57888
rect 63957 57879 64015 57885
rect 64601 57885 64613 57888
rect 64647 57885 64659 57919
rect 64601 57879 64659 57885
rect 64049 57783 64107 57789
rect 64049 57749 64061 57783
rect 64095 57780 64107 57783
rect 64230 57780 64236 57792
rect 64095 57752 64236 57780
rect 64095 57749 64107 57752
rect 64049 57743 64107 57749
rect 64230 57740 64236 57752
rect 64288 57740 64294 57792
rect 1104 57690 68816 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 68816 57690
rect 1104 57616 68816 57638
rect 34698 57508 34704 57520
rect 34256 57480 34704 57508
rect 34256 57449 34284 57480
rect 34698 57468 34704 57480
rect 34756 57468 34762 57520
rect 64230 57508 64236 57520
rect 64191 57480 64236 57508
rect 64230 57468 64236 57480
rect 64288 57468 64294 57520
rect 65889 57511 65947 57517
rect 65889 57477 65901 57511
rect 65935 57508 65947 57511
rect 66162 57508 66168 57520
rect 65935 57480 66168 57508
rect 65935 57477 65947 57480
rect 65889 57471 65947 57477
rect 66162 57468 66168 57480
rect 66220 57468 66226 57520
rect 34241 57443 34299 57449
rect 34241 57409 34253 57443
rect 34287 57409 34299 57443
rect 34241 57403 34299 57409
rect 63494 57400 63500 57452
rect 63552 57440 63558 57452
rect 64049 57443 64107 57449
rect 64049 57440 64061 57443
rect 63552 57412 64061 57440
rect 63552 57400 63558 57412
rect 64049 57409 64061 57412
rect 64095 57409 64107 57443
rect 64049 57403 64107 57409
rect 34422 57372 34428 57384
rect 34383 57344 34428 57372
rect 34422 57332 34428 57344
rect 34480 57332 34486 57384
rect 35802 57372 35808 57384
rect 35763 57344 35808 57372
rect 35802 57332 35808 57344
rect 35860 57332 35866 57384
rect 1104 57146 68816 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 68816 57146
rect 1104 57072 68816 57094
rect 34422 56992 34428 57044
rect 34480 57032 34486 57044
rect 34793 57035 34851 57041
rect 34793 57032 34805 57035
rect 34480 57004 34805 57032
rect 34480 56992 34486 57004
rect 34793 57001 34805 57004
rect 34839 57001 34851 57035
rect 34793 56995 34851 57001
rect 34885 56831 34943 56837
rect 34885 56797 34897 56831
rect 34931 56828 34943 56831
rect 35434 56828 35440 56840
rect 34931 56800 35440 56828
rect 34931 56797 34943 56800
rect 34885 56791 34943 56797
rect 35434 56788 35440 56800
rect 35492 56788 35498 56840
rect 49234 56828 49240 56840
rect 49195 56800 49240 56828
rect 49234 56788 49240 56800
rect 49292 56788 49298 56840
rect 63954 56788 63960 56840
rect 64012 56828 64018 56840
rect 64049 56831 64107 56837
rect 64049 56828 64061 56831
rect 64012 56800 64061 56828
rect 64012 56788 64018 56800
rect 64049 56797 64061 56800
rect 64095 56797 64107 56831
rect 64049 56791 64107 56797
rect 1104 56602 68816 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 68816 56602
rect 1104 56528 68816 56550
rect 63586 56448 63592 56500
rect 63644 56488 63650 56500
rect 64414 56488 64420 56500
rect 63644 56460 64420 56488
rect 63644 56448 63650 56460
rect 64414 56448 64420 56460
rect 64472 56448 64478 56500
rect 49234 56352 49240 56364
rect 49195 56324 49240 56352
rect 49234 56312 49240 56324
rect 49292 56312 49298 56364
rect 63954 56352 63960 56364
rect 63915 56324 63960 56352
rect 63954 56312 63960 56324
rect 64012 56312 64018 56364
rect 2774 56244 2780 56296
rect 2832 56284 2838 56296
rect 32950 56284 32956 56296
rect 2832 56256 26234 56284
rect 32911 56256 32956 56284
rect 2832 56244 2838 56256
rect 26206 56216 26234 56256
rect 32950 56244 32956 56256
rect 33008 56244 33014 56296
rect 33134 56284 33140 56296
rect 33095 56256 33140 56284
rect 33134 56244 33140 56256
rect 33192 56244 33198 56296
rect 33413 56287 33471 56293
rect 33413 56253 33425 56287
rect 33459 56253 33471 56287
rect 33413 56247 33471 56253
rect 49421 56287 49479 56293
rect 49421 56253 49433 56287
rect 49467 56253 49479 56287
rect 49421 56247 49479 56253
rect 51077 56287 51135 56293
rect 51077 56253 51089 56287
rect 51123 56284 51135 56287
rect 64141 56287 64199 56293
rect 51123 56256 55214 56284
rect 51123 56253 51135 56256
rect 51077 56247 51135 56253
rect 33428 56216 33456 56247
rect 26206 56188 33456 56216
rect 49234 56176 49240 56228
rect 49292 56216 49298 56228
rect 49436 56216 49464 56247
rect 49292 56188 49464 56216
rect 55186 56216 55214 56256
rect 64141 56253 64153 56287
rect 64187 56284 64199 56287
rect 64230 56284 64236 56296
rect 64187 56256 64236 56284
rect 64187 56253 64199 56256
rect 64141 56247 64199 56253
rect 64230 56244 64236 56256
rect 64288 56244 64294 56296
rect 64414 56284 64420 56296
rect 64375 56256 64420 56284
rect 64414 56244 64420 56256
rect 64472 56244 64478 56296
rect 66162 56216 66168 56228
rect 55186 56188 66168 56216
rect 49292 56176 49298 56188
rect 66162 56176 66168 56188
rect 66220 56176 66226 56228
rect 1104 56058 68816 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 68816 56058
rect 1104 55984 68816 56006
rect 32950 55944 32956 55956
rect 32911 55916 32956 55944
rect 32950 55904 32956 55916
rect 33008 55904 33014 55956
rect 49234 55944 49240 55956
rect 49195 55916 49240 55944
rect 49234 55904 49240 55916
rect 49292 55904 49298 55956
rect 64230 55944 64236 55956
rect 64191 55916 64236 55944
rect 64230 55904 64236 55916
rect 64288 55904 64294 55956
rect 45526 55780 49188 55808
rect 33781 55743 33839 55749
rect 33781 55709 33793 55743
rect 33827 55740 33839 55743
rect 35342 55740 35348 55752
rect 33827 55712 35348 55740
rect 33827 55709 33839 55712
rect 33781 55703 33839 55709
rect 35342 55700 35348 55712
rect 35400 55700 35406 55752
rect 35434 55700 35440 55752
rect 35492 55740 35498 55752
rect 45526 55740 45554 55780
rect 48682 55740 48688 55752
rect 35492 55712 45554 55740
rect 48643 55712 48688 55740
rect 35492 55700 35498 55712
rect 48682 55700 48688 55712
rect 48740 55700 48746 55752
rect 49160 55749 49188 55780
rect 49145 55743 49203 55749
rect 49145 55709 49157 55743
rect 49191 55709 49203 55743
rect 63678 55740 63684 55752
rect 63639 55712 63684 55740
rect 49145 55703 49203 55709
rect 63678 55700 63684 55712
rect 63736 55700 63742 55752
rect 64325 55743 64383 55749
rect 64325 55709 64337 55743
rect 64371 55740 64383 55743
rect 64690 55740 64696 55752
rect 64371 55712 64696 55740
rect 64371 55709 64383 55712
rect 64325 55703 64383 55709
rect 64690 55700 64696 55712
rect 64748 55740 64754 55752
rect 64877 55743 64935 55749
rect 64877 55740 64889 55743
rect 64748 55712 64889 55740
rect 64748 55700 64754 55712
rect 64877 55709 64889 55712
rect 64923 55709 64935 55743
rect 64877 55703 64935 55709
rect 64966 55700 64972 55752
rect 65024 55740 65030 55752
rect 65613 55743 65671 55749
rect 65613 55740 65625 55743
rect 65024 55712 65625 55740
rect 65024 55700 65030 55712
rect 65613 55709 65625 55712
rect 65659 55709 65671 55743
rect 65613 55703 65671 55709
rect 63586 55604 63592 55616
rect 63547 55576 63592 55604
rect 63586 55564 63592 55576
rect 63644 55564 63650 55616
rect 64969 55607 65027 55613
rect 64969 55573 64981 55607
rect 65015 55604 65027 55607
rect 65150 55604 65156 55616
rect 65015 55576 65156 55604
rect 65015 55573 65027 55576
rect 64969 55567 65027 55573
rect 65150 55564 65156 55576
rect 65208 55564 65214 55616
rect 1104 55514 68816 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 68816 55514
rect 1104 55440 68816 55462
rect 50525 55335 50583 55341
rect 50525 55301 50537 55335
rect 50571 55332 50583 55335
rect 50614 55332 50620 55344
rect 50571 55304 50620 55332
rect 50571 55301 50583 55304
rect 50525 55295 50583 55301
rect 50614 55292 50620 55304
rect 50672 55292 50678 55344
rect 65150 55332 65156 55344
rect 65111 55304 65156 55332
rect 65150 55292 65156 55304
rect 65208 55292 65214 55344
rect 66806 55332 66812 55344
rect 66767 55304 66812 55332
rect 66806 55292 66812 55304
rect 66864 55292 66870 55344
rect 3326 55224 3332 55276
rect 3384 55264 3390 55276
rect 33505 55267 33563 55273
rect 33505 55264 33517 55267
rect 3384 55236 33517 55264
rect 3384 55224 3390 55236
rect 33505 55233 33517 55236
rect 33551 55233 33563 55267
rect 33505 55227 33563 55233
rect 35342 55224 35348 55276
rect 35400 55264 35406 55276
rect 48682 55264 48688 55276
rect 35400 55236 35445 55264
rect 48643 55236 48688 55264
rect 35400 55224 35406 55236
rect 48682 55224 48688 55236
rect 48740 55224 48746 55276
rect 64966 55264 64972 55276
rect 64927 55236 64972 55264
rect 64966 55224 64972 55236
rect 65024 55224 65030 55276
rect 34790 55156 34796 55208
rect 34848 55196 34854 55208
rect 35161 55199 35219 55205
rect 35161 55196 35173 55199
rect 34848 55168 35173 55196
rect 34848 55156 34854 55168
rect 35161 55165 35173 55168
rect 35207 55165 35219 55199
rect 48866 55196 48872 55208
rect 48827 55168 48872 55196
rect 35161 55159 35219 55165
rect 48866 55156 48872 55168
rect 48924 55156 48930 55208
rect 63218 55020 63224 55072
rect 63276 55060 63282 55072
rect 63681 55063 63739 55069
rect 63681 55060 63693 55063
rect 63276 55032 63693 55060
rect 63276 55020 63282 55032
rect 63681 55029 63693 55032
rect 63727 55029 63739 55063
rect 63681 55023 63739 55029
rect 1104 54970 68816 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 68816 54970
rect 1104 54896 68816 54918
rect 33134 54816 33140 54868
rect 33192 54856 33198 54868
rect 33597 54859 33655 54865
rect 33597 54856 33609 54859
rect 33192 54828 33609 54856
rect 33192 54816 33198 54828
rect 33597 54825 33609 54828
rect 33643 54825 33655 54859
rect 34790 54856 34796 54868
rect 34751 54828 34796 54856
rect 33597 54819 33655 54825
rect 34790 54816 34796 54828
rect 34848 54816 34854 54868
rect 48685 54859 48743 54865
rect 48685 54825 48697 54859
rect 48731 54856 48743 54859
rect 48866 54856 48872 54868
rect 48731 54828 48872 54856
rect 48731 54825 48743 54828
rect 48685 54819 48743 54825
rect 48866 54816 48872 54828
rect 48924 54816 48930 54868
rect 63218 54720 63224 54732
rect 63179 54692 63224 54720
rect 63218 54680 63224 54692
rect 63276 54680 63282 54732
rect 63405 54723 63463 54729
rect 63405 54689 63417 54723
rect 63451 54720 63463 54723
rect 63586 54720 63592 54732
rect 63451 54692 63592 54720
rect 63451 54689 63463 54692
rect 63405 54683 63463 54689
rect 63586 54680 63592 54692
rect 63644 54680 63650 54732
rect 65058 54720 65064 54732
rect 65019 54692 65064 54720
rect 65058 54680 65064 54692
rect 65116 54680 65122 54732
rect 33689 54655 33747 54661
rect 33689 54621 33701 54655
rect 33735 54621 33747 54655
rect 33689 54615 33747 54621
rect 34885 54655 34943 54661
rect 34885 54621 34897 54655
rect 34931 54652 34943 54655
rect 38010 54652 38016 54664
rect 34931 54624 38016 54652
rect 34931 54621 34943 54624
rect 34885 54615 34943 54621
rect 33704 54584 33732 54615
rect 38010 54612 38016 54624
rect 38068 54612 38074 54664
rect 48590 54652 48596 54664
rect 48551 54624 48596 54652
rect 48590 54612 48596 54624
rect 48648 54612 48654 54664
rect 40770 54584 40776 54596
rect 33704 54556 40776 54584
rect 40770 54544 40776 54556
rect 40828 54544 40834 54596
rect 1104 54426 68816 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 68816 54426
rect 1104 54352 68816 54374
rect 1104 53882 68816 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 68816 53882
rect 1104 53808 68816 53830
rect 1104 53338 68816 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 68816 53338
rect 1104 53264 68816 53286
rect 40678 52844 40684 52896
rect 40736 52884 40742 52896
rect 40773 52887 40831 52893
rect 40773 52884 40785 52887
rect 40736 52856 40785 52884
rect 40736 52844 40742 52856
rect 40773 52853 40785 52856
rect 40819 52853 40831 52887
rect 40773 52847 40831 52853
rect 1104 52794 68816 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 68816 52794
rect 1104 52720 68816 52742
rect 40126 52572 40132 52624
rect 40184 52612 40190 52624
rect 40184 52584 41184 52612
rect 40184 52572 40190 52584
rect 40678 52544 40684 52556
rect 40639 52516 40684 52544
rect 40678 52504 40684 52516
rect 40736 52504 40742 52556
rect 41156 52553 41184 52584
rect 41141 52547 41199 52553
rect 41141 52513 41153 52547
rect 41187 52513 41199 52547
rect 41141 52507 41199 52513
rect 40862 52408 40868 52420
rect 40823 52380 40868 52408
rect 40862 52368 40868 52380
rect 40920 52368 40926 52420
rect 1104 52250 68816 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 68816 52250
rect 1104 52176 68816 52198
rect 40862 52136 40868 52148
rect 40823 52108 40868 52136
rect 40862 52096 40868 52108
rect 40920 52096 40926 52148
rect 40770 52000 40776 52012
rect 40731 51972 40776 52000
rect 40770 51960 40776 51972
rect 40828 51960 40834 52012
rect 31573 51935 31631 51941
rect 31573 51901 31585 51935
rect 31619 51932 31631 51935
rect 32125 51935 32183 51941
rect 32125 51932 32137 51935
rect 31619 51904 32137 51932
rect 31619 51901 31631 51904
rect 31573 51895 31631 51901
rect 32125 51901 32137 51904
rect 32171 51901 32183 51935
rect 32306 51932 32312 51944
rect 32267 51904 32312 51932
rect 32125 51895 32183 51901
rect 32306 51892 32312 51904
rect 32364 51892 32370 51944
rect 32585 51935 32643 51941
rect 32585 51901 32597 51935
rect 32631 51901 32643 51935
rect 32585 51895 32643 51901
rect 31754 51824 31760 51876
rect 31812 51864 31818 51876
rect 32600 51864 32628 51895
rect 31812 51836 32628 51864
rect 31812 51824 31818 51836
rect 50982 51756 50988 51808
rect 51040 51796 51046 51808
rect 51077 51799 51135 51805
rect 51077 51796 51089 51799
rect 51040 51768 51089 51796
rect 51040 51756 51046 51768
rect 51077 51765 51089 51768
rect 51123 51765 51135 51799
rect 51077 51759 51135 51765
rect 1104 51706 68816 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 68816 51706
rect 1104 51632 68816 51654
rect 31849 51595 31907 51601
rect 31849 51561 31861 51595
rect 31895 51592 31907 51595
rect 32306 51592 32312 51604
rect 31895 51564 32312 51592
rect 31895 51561 31907 51564
rect 31849 51555 31907 51561
rect 32306 51552 32312 51564
rect 32364 51552 32370 51604
rect 50982 51456 50988 51468
rect 50943 51428 50988 51456
rect 50982 51416 50988 51428
rect 51040 51416 51046 51468
rect 52822 51456 52828 51468
rect 52783 51428 52828 51456
rect 52822 51416 52828 51428
rect 52880 51416 52886 51468
rect 31757 51391 31815 51397
rect 31757 51357 31769 51391
rect 31803 51388 31815 51391
rect 31803 51360 35894 51388
rect 31803 51357 31815 51360
rect 31757 51351 31815 51357
rect 35866 51252 35894 51360
rect 51166 51320 51172 51332
rect 51127 51292 51172 51320
rect 51166 51280 51172 51292
rect 51224 51280 51230 51332
rect 37918 51252 37924 51264
rect 35866 51224 37924 51252
rect 37918 51212 37924 51224
rect 37976 51252 37982 51264
rect 48590 51252 48596 51264
rect 37976 51224 48596 51252
rect 37976 51212 37982 51224
rect 48590 51212 48596 51224
rect 48648 51252 48654 51264
rect 48958 51252 48964 51264
rect 48648 51224 48964 51252
rect 48648 51212 48654 51224
rect 48958 51212 48964 51224
rect 49016 51212 49022 51264
rect 1104 51162 68816 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 68816 51162
rect 1104 51088 68816 51110
rect 50801 51051 50859 51057
rect 50801 51017 50813 51051
rect 50847 51048 50859 51051
rect 51166 51048 51172 51060
rect 50847 51020 51172 51048
rect 50847 51017 50859 51020
rect 50801 51011 50859 51017
rect 51166 51008 51172 51020
rect 51224 51008 51230 51060
rect 43438 50872 43444 50924
rect 43496 50912 43502 50924
rect 50709 50915 50767 50921
rect 50709 50912 50721 50915
rect 43496 50884 50721 50912
rect 43496 50872 43502 50884
rect 50709 50881 50721 50884
rect 50755 50881 50767 50915
rect 50709 50875 50767 50881
rect 24394 50668 24400 50720
rect 24452 50708 24458 50720
rect 24489 50711 24547 50717
rect 24489 50708 24501 50711
rect 24452 50680 24501 50708
rect 24452 50668 24458 50680
rect 24489 50677 24501 50680
rect 24535 50677 24547 50711
rect 24489 50671 24547 50677
rect 1104 50618 68816 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 68816 50618
rect 1104 50544 68816 50566
rect 6914 50328 6920 50380
rect 6972 50368 6978 50380
rect 24857 50371 24915 50377
rect 24857 50368 24869 50371
rect 6972 50340 24869 50368
rect 6972 50328 6978 50340
rect 24857 50337 24869 50340
rect 24903 50337 24915 50371
rect 24857 50331 24915 50337
rect 24394 50300 24400 50312
rect 24355 50272 24400 50300
rect 24394 50260 24400 50272
rect 24452 50260 24458 50312
rect 24581 50235 24639 50241
rect 24581 50201 24593 50235
rect 24627 50232 24639 50235
rect 24854 50232 24860 50244
rect 24627 50204 24860 50232
rect 24627 50201 24639 50204
rect 24581 50195 24639 50201
rect 24854 50192 24860 50204
rect 24912 50192 24918 50244
rect 1104 50074 68816 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 68816 50074
rect 1104 50000 68816 50022
rect 24854 49960 24860 49972
rect 24815 49932 24860 49960
rect 24854 49920 24860 49932
rect 24912 49920 24918 49972
rect 24949 49827 25007 49833
rect 24949 49793 24961 49827
rect 24995 49824 25007 49827
rect 35342 49824 35348 49836
rect 24995 49796 35348 49824
rect 24995 49793 25007 49796
rect 24949 49787 25007 49793
rect 35342 49784 35348 49796
rect 35400 49784 35406 49836
rect 1104 49530 68816 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 68816 49530
rect 1104 49456 68816 49478
rect 54110 49172 54116 49224
rect 54168 49212 54174 49224
rect 54205 49215 54263 49221
rect 54205 49212 54217 49215
rect 54168 49184 54217 49212
rect 54168 49172 54174 49184
rect 54205 49181 54217 49184
rect 54251 49181 54263 49215
rect 54205 49175 54263 49181
rect 1104 48986 68816 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 68816 48986
rect 1104 48912 68816 48934
rect 51074 48696 51080 48748
rect 51132 48736 51138 48748
rect 53469 48739 53527 48745
rect 53469 48736 53481 48739
rect 51132 48708 53481 48736
rect 51132 48696 51138 48708
rect 53469 48705 53481 48708
rect 53515 48705 53527 48739
rect 54110 48736 54116 48748
rect 54071 48708 54116 48736
rect 53469 48699 53527 48705
rect 54110 48696 54116 48708
rect 54168 48696 54174 48748
rect 53561 48671 53619 48677
rect 53561 48637 53573 48671
rect 53607 48668 53619 48671
rect 54297 48671 54355 48677
rect 54297 48668 54309 48671
rect 53607 48640 54309 48668
rect 53607 48637 53619 48640
rect 53561 48631 53619 48637
rect 54297 48637 54309 48640
rect 54343 48637 54355 48671
rect 54297 48631 54355 48637
rect 55953 48671 56011 48677
rect 55953 48637 55965 48671
rect 55999 48668 56011 48671
rect 65426 48668 65432 48680
rect 55999 48640 65432 48668
rect 55999 48637 56011 48640
rect 55953 48631 56011 48637
rect 65426 48628 65432 48640
rect 65484 48628 65490 48680
rect 20993 48535 21051 48541
rect 20993 48501 21005 48535
rect 21039 48532 21051 48535
rect 22646 48532 22652 48544
rect 21039 48504 22652 48532
rect 21039 48501 21051 48504
rect 20993 48495 21051 48501
rect 22646 48492 22652 48504
rect 22704 48492 22710 48544
rect 1104 48442 68816 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 68816 48442
rect 1104 48368 68816 48390
rect 22646 48192 22652 48204
rect 22607 48164 22652 48192
rect 22646 48152 22652 48164
rect 22704 48152 22710 48204
rect 3694 48016 3700 48068
rect 3752 48056 3758 48068
rect 20809 48059 20867 48065
rect 20809 48056 20821 48059
rect 3752 48028 20821 48056
rect 3752 48016 3758 48028
rect 20809 48025 20821 48028
rect 20855 48025 20867 48059
rect 20809 48019 20867 48025
rect 21910 48016 21916 48068
rect 21968 48056 21974 48068
rect 22465 48059 22523 48065
rect 22465 48056 22477 48059
rect 21968 48028 22477 48056
rect 21968 48016 21974 48028
rect 22465 48025 22477 48028
rect 22511 48025 22523 48059
rect 22465 48019 22523 48025
rect 1104 47898 68816 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 68816 47898
rect 1104 47824 68816 47846
rect 21910 47784 21916 47796
rect 21871 47756 21916 47784
rect 21910 47744 21916 47756
rect 21968 47744 21974 47796
rect 49418 47716 49424 47728
rect 49379 47688 49424 47716
rect 49418 47676 49424 47688
rect 49476 47676 49482 47728
rect 22002 47648 22008 47660
rect 21963 47620 22008 47648
rect 22002 47608 22008 47620
rect 22060 47608 22066 47660
rect 47029 47583 47087 47589
rect 47029 47549 47041 47583
rect 47075 47580 47087 47583
rect 47581 47583 47639 47589
rect 47581 47580 47593 47583
rect 47075 47552 47593 47580
rect 47075 47549 47087 47552
rect 47029 47543 47087 47549
rect 47581 47549 47593 47552
rect 47627 47549 47639 47583
rect 47762 47580 47768 47592
rect 47723 47552 47768 47580
rect 47581 47543 47639 47549
rect 47762 47540 47768 47552
rect 47820 47540 47826 47592
rect 61930 47444 61936 47456
rect 61891 47416 61936 47444
rect 61930 47404 61936 47416
rect 61988 47404 61994 47456
rect 1104 47354 68816 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 68816 47354
rect 1104 47280 68816 47302
rect 46937 47243 46995 47249
rect 46937 47209 46949 47243
rect 46983 47240 46995 47243
rect 47762 47240 47768 47252
rect 46983 47212 47768 47240
rect 46983 47209 46995 47212
rect 46937 47203 46995 47209
rect 47762 47200 47768 47212
rect 47820 47200 47826 47252
rect 66162 47172 66168 47184
rect 59740 47144 66168 47172
rect 57885 47107 57943 47113
rect 57885 47073 57897 47107
rect 57931 47104 57943 47107
rect 58066 47104 58072 47116
rect 57931 47076 58072 47104
rect 57931 47073 57943 47076
rect 57885 47067 57943 47073
rect 58066 47064 58072 47076
rect 58124 47064 58130 47116
rect 59740 47113 59768 47144
rect 66162 47132 66168 47144
rect 66220 47132 66226 47184
rect 59725 47107 59783 47113
rect 59725 47073 59737 47107
rect 59771 47073 59783 47107
rect 61930 47104 61936 47116
rect 61891 47076 61936 47104
rect 59725 47067 59783 47073
rect 61930 47064 61936 47076
rect 61988 47064 61994 47116
rect 63773 47107 63831 47113
rect 63773 47073 63785 47107
rect 63819 47104 63831 47107
rect 64782 47104 64788 47116
rect 63819 47076 64788 47104
rect 63819 47073 63831 47076
rect 63773 47067 63831 47073
rect 64782 47064 64788 47076
rect 64840 47064 64846 47116
rect 44910 46996 44916 47048
rect 44968 47036 44974 47048
rect 46845 47039 46903 47045
rect 46845 47036 46857 47039
rect 44968 47008 46857 47036
rect 44968 46996 44974 47008
rect 46845 47005 46857 47008
rect 46891 47005 46903 47039
rect 56502 47036 56508 47048
rect 46845 46999 46903 47005
rect 55186 47008 56508 47036
rect 40770 46928 40776 46980
rect 40828 46968 40834 46980
rect 55186 46968 55214 47008
rect 56502 46996 56508 47008
rect 56560 47036 56566 47048
rect 57241 47039 57299 47045
rect 57241 47036 57253 47039
rect 56560 47008 57253 47036
rect 56560 46996 56566 47008
rect 57241 47005 57253 47008
rect 57287 47005 57299 47039
rect 57241 46999 57299 47005
rect 40828 46940 55214 46968
rect 57333 46971 57391 46977
rect 40828 46928 40834 46940
rect 57333 46937 57345 46971
rect 57379 46968 57391 46971
rect 58069 46971 58127 46977
rect 58069 46968 58081 46971
rect 57379 46940 58081 46968
rect 57379 46937 57391 46940
rect 57333 46931 57391 46937
rect 58069 46937 58081 46940
rect 58115 46937 58127 46971
rect 62114 46968 62120 46980
rect 62075 46940 62120 46968
rect 58069 46931 58127 46937
rect 62114 46928 62120 46940
rect 62172 46928 62178 46980
rect 1104 46810 68816 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 68816 46810
rect 1104 46736 68816 46758
rect 61749 46699 61807 46705
rect 61749 46665 61761 46699
rect 61795 46696 61807 46699
rect 62114 46696 62120 46708
rect 61795 46668 62120 46696
rect 61795 46665 61807 46668
rect 61749 46659 61807 46665
rect 62114 46656 62120 46668
rect 62172 46656 62178 46708
rect 57977 46563 58035 46569
rect 57977 46529 57989 46563
rect 58023 46560 58035 46563
rect 58066 46560 58072 46572
rect 58023 46532 58072 46560
rect 58023 46529 58035 46532
rect 57977 46523 58035 46529
rect 58066 46520 58072 46532
rect 58124 46520 58130 46572
rect 60918 46520 60924 46572
rect 60976 46560 60982 46572
rect 61657 46563 61715 46569
rect 61657 46560 61669 46563
rect 60976 46532 61669 46560
rect 60976 46520 60982 46532
rect 61657 46529 61669 46532
rect 61703 46529 61715 46563
rect 61657 46523 61715 46529
rect 41414 46452 41420 46504
rect 41472 46492 41478 46504
rect 42426 46492 42432 46504
rect 41472 46464 42432 46492
rect 41472 46452 41478 46464
rect 42426 46452 42432 46464
rect 42484 46452 42490 46504
rect 41966 46316 41972 46368
rect 42024 46356 42030 46368
rect 42429 46359 42487 46365
rect 42429 46356 42441 46359
rect 42024 46328 42441 46356
rect 42024 46316 42030 46328
rect 42429 46325 42441 46328
rect 42475 46325 42487 46359
rect 42429 46319 42487 46325
rect 1104 46266 68816 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 68816 46266
rect 1104 46192 68816 46214
rect 51074 46084 51080 46096
rect 41340 46056 51080 46084
rect 35526 45908 35532 45960
rect 35584 45948 35590 45960
rect 41340 45957 41368 46056
rect 51074 46044 51080 46056
rect 51132 46044 51138 46096
rect 41966 46016 41972 46028
rect 41927 45988 41972 46016
rect 41966 45976 41972 45988
rect 42024 45976 42030 46028
rect 42426 46016 42432 46028
rect 42387 45988 42432 46016
rect 42426 45976 42432 45988
rect 42484 45976 42490 46028
rect 41325 45951 41383 45957
rect 41325 45948 41337 45951
rect 35584 45920 41337 45948
rect 35584 45908 35590 45920
rect 41325 45917 41337 45920
rect 41371 45917 41383 45951
rect 61010 45948 61016 45960
rect 60971 45920 61016 45948
rect 41325 45911 41383 45917
rect 61010 45908 61016 45920
rect 61068 45908 61074 45960
rect 41417 45883 41475 45889
rect 41417 45849 41429 45883
rect 41463 45880 41475 45883
rect 42153 45883 42211 45889
rect 42153 45880 42165 45883
rect 41463 45852 42165 45880
rect 41463 45849 41475 45852
rect 41417 45843 41475 45849
rect 42153 45849 42165 45852
rect 42199 45849 42211 45883
rect 42153 45843 42211 45849
rect 1104 45722 68816 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 68816 45722
rect 1104 45648 68816 45670
rect 61010 45540 61016 45552
rect 60660 45512 61016 45540
rect 60660 45481 60688 45512
rect 61010 45500 61016 45512
rect 61068 45500 61074 45552
rect 62485 45543 62543 45549
rect 62485 45509 62497 45543
rect 62531 45540 62543 45543
rect 65978 45540 65984 45552
rect 62531 45512 65984 45540
rect 62531 45509 62543 45512
rect 62485 45503 62543 45509
rect 65978 45500 65984 45512
rect 66036 45500 66042 45552
rect 60645 45475 60703 45481
rect 60645 45441 60657 45475
rect 60691 45441 60703 45475
rect 60645 45435 60703 45441
rect 60826 45404 60832 45416
rect 60787 45376 60832 45404
rect 60826 45364 60832 45376
rect 60884 45364 60890 45416
rect 1104 45178 68816 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 68816 45178
rect 1104 45104 68816 45126
rect 60645 45067 60703 45073
rect 60645 45033 60657 45067
rect 60691 45064 60703 45067
rect 60826 45064 60832 45076
rect 60691 45036 60832 45064
rect 60691 45033 60703 45036
rect 60645 45027 60703 45033
rect 60826 45024 60832 45036
rect 60884 45024 60890 45076
rect 60550 44860 60556 44872
rect 60511 44832 60556 44860
rect 60550 44820 60556 44832
rect 60608 44820 60614 44872
rect 1104 44634 68816 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 68816 44634
rect 1104 44560 68816 44582
rect 1104 44090 68816 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 68816 44090
rect 1104 44016 68816 44038
rect 60274 43732 60280 43784
rect 60332 43772 60338 43784
rect 60461 43775 60519 43781
rect 60461 43772 60473 43775
rect 60332 43744 60473 43772
rect 60332 43732 60338 43744
rect 60461 43741 60473 43744
rect 60507 43741 60519 43775
rect 60461 43735 60519 43741
rect 1104 43546 68816 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 68816 43546
rect 1104 43472 68816 43494
rect 60274 43296 60280 43308
rect 60235 43268 60280 43296
rect 60274 43256 60280 43268
rect 60332 43256 60338 43308
rect 60458 43228 60464 43240
rect 60419 43200 60464 43228
rect 60458 43188 60464 43200
rect 60516 43188 60522 43240
rect 62022 43228 62028 43240
rect 61983 43200 62028 43228
rect 62022 43188 62028 43200
rect 62080 43188 62086 43240
rect 16758 43052 16764 43104
rect 16816 43092 16822 43104
rect 16853 43095 16911 43101
rect 16853 43092 16865 43095
rect 16816 43064 16865 43092
rect 16816 43052 16822 43064
rect 16853 43061 16865 43064
rect 16899 43061 16911 43095
rect 16853 43055 16911 43061
rect 34149 43095 34207 43101
rect 34149 43061 34161 43095
rect 34195 43092 34207 43095
rect 34698 43092 34704 43104
rect 34195 43064 34704 43092
rect 34195 43061 34207 43064
rect 34149 43055 34207 43061
rect 34698 43052 34704 43064
rect 34756 43052 34762 43104
rect 45002 43052 45008 43104
rect 45060 43092 45066 43104
rect 45097 43095 45155 43101
rect 45097 43092 45109 43095
rect 45060 43064 45109 43092
rect 45060 43052 45066 43064
rect 45097 43061 45109 43064
rect 45143 43061 45155 43095
rect 52730 43092 52736 43104
rect 52691 43064 52736 43092
rect 45097 43055 45155 43061
rect 52730 43052 52736 43064
rect 52788 43052 52794 43104
rect 1104 43002 68816 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 68816 43002
rect 1104 42928 68816 42950
rect 60458 42848 60464 42900
rect 60516 42888 60522 42900
rect 60553 42891 60611 42897
rect 60553 42888 60565 42891
rect 60516 42860 60565 42888
rect 60516 42848 60522 42860
rect 60553 42857 60565 42860
rect 60599 42857 60611 42891
rect 60553 42851 60611 42857
rect 3694 42712 3700 42764
rect 3752 42752 3758 42764
rect 35161 42755 35219 42761
rect 35161 42752 35173 42755
rect 3752 42724 35173 42752
rect 3752 42712 3758 42724
rect 35161 42721 35173 42724
rect 35207 42721 35219 42755
rect 45002 42752 45008 42764
rect 44963 42724 45008 42752
rect 35161 42715 35219 42721
rect 45002 42712 45008 42724
rect 45060 42712 45066 42764
rect 46842 42752 46848 42764
rect 46803 42724 46848 42752
rect 46842 42712 46848 42724
rect 46900 42712 46906 42764
rect 52181 42755 52239 42761
rect 52181 42721 52193 42755
rect 52227 42752 52239 42755
rect 52730 42752 52736 42764
rect 52227 42724 52736 42752
rect 52227 42721 52239 42724
rect 52181 42715 52239 42721
rect 52730 42712 52736 42724
rect 52788 42712 52794 42764
rect 16758 42684 16764 42696
rect 16719 42656 16764 42684
rect 16758 42644 16764 42656
rect 16816 42644 16822 42696
rect 34698 42684 34704 42696
rect 34659 42656 34704 42684
rect 34698 42644 34704 42656
rect 34756 42644 34762 42696
rect 48958 42644 48964 42696
rect 49016 42684 49022 42696
rect 51537 42687 51595 42693
rect 51537 42684 51549 42687
rect 49016 42656 51549 42684
rect 49016 42644 49022 42656
rect 51537 42653 51549 42656
rect 51583 42653 51595 42687
rect 51537 42647 51595 42653
rect 59722 42644 59728 42696
rect 59780 42684 59786 42696
rect 60461 42687 60519 42693
rect 60461 42684 60473 42687
rect 59780 42656 60473 42684
rect 59780 42644 59786 42656
rect 60461 42653 60473 42656
rect 60507 42684 60519 42687
rect 60550 42684 60556 42696
rect 60507 42656 60556 42684
rect 60507 42653 60519 42656
rect 60461 42647 60519 42653
rect 60550 42644 60556 42656
rect 60608 42644 60614 42696
rect 16942 42616 16948 42628
rect 16903 42588 16948 42616
rect 16942 42576 16948 42588
rect 17000 42576 17006 42628
rect 18601 42619 18659 42625
rect 18601 42585 18613 42619
rect 18647 42585 18659 42619
rect 18601 42579 18659 42585
rect 16574 42508 16580 42560
rect 16632 42548 16638 42560
rect 18616 42548 18644 42579
rect 34606 42576 34612 42628
rect 34664 42616 34670 42628
rect 34885 42619 34943 42625
rect 34885 42616 34897 42619
rect 34664 42588 34897 42616
rect 34664 42576 34670 42588
rect 34885 42585 34897 42588
rect 34931 42585 34943 42619
rect 34885 42579 34943 42585
rect 45002 42576 45008 42628
rect 45060 42616 45066 42628
rect 45189 42619 45247 42625
rect 45189 42616 45201 42619
rect 45060 42588 45201 42616
rect 45060 42576 45066 42588
rect 45189 42585 45201 42588
rect 45235 42585 45247 42619
rect 45189 42579 45247 42585
rect 51629 42619 51687 42625
rect 51629 42585 51641 42619
rect 51675 42616 51687 42619
rect 52365 42619 52423 42625
rect 52365 42616 52377 42619
rect 51675 42588 52377 42616
rect 51675 42585 51687 42588
rect 51629 42579 51687 42585
rect 52365 42585 52377 42588
rect 52411 42585 52423 42619
rect 52365 42579 52423 42585
rect 54021 42619 54079 42625
rect 54021 42585 54033 42619
rect 54067 42616 54079 42619
rect 66162 42616 66168 42628
rect 54067 42588 66168 42616
rect 54067 42585 54079 42588
rect 54021 42579 54079 42585
rect 66162 42576 66168 42588
rect 66220 42576 66226 42628
rect 16632 42520 18644 42548
rect 16632 42508 16638 42520
rect 1104 42458 68816 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 68816 42458
rect 1104 42384 68816 42406
rect 16942 42344 16948 42356
rect 16903 42316 16948 42344
rect 16942 42304 16948 42316
rect 17000 42304 17006 42356
rect 34606 42344 34612 42356
rect 34567 42316 34612 42344
rect 34606 42304 34612 42316
rect 34664 42304 34670 42356
rect 45002 42344 45008 42356
rect 44963 42316 45008 42344
rect 45002 42304 45008 42316
rect 45060 42304 45066 42356
rect 14458 42168 14464 42220
rect 14516 42208 14522 42220
rect 16853 42211 16911 42217
rect 16853 42208 16865 42211
rect 14516 42180 16865 42208
rect 14516 42168 14522 42180
rect 16853 42177 16865 42180
rect 16899 42208 16911 42211
rect 32858 42208 32864 42220
rect 16899 42180 32864 42208
rect 16899 42177 16911 42180
rect 16853 42171 16911 42177
rect 32858 42168 32864 42180
rect 32916 42168 32922 42220
rect 34701 42211 34759 42217
rect 34701 42177 34713 42211
rect 34747 42208 34759 42211
rect 34747 42180 35894 42208
rect 34747 42177 34759 42180
rect 34701 42171 34759 42177
rect 35866 42140 35894 42180
rect 38194 42168 38200 42220
rect 38252 42208 38258 42220
rect 44910 42208 44916 42220
rect 38252 42180 44916 42208
rect 38252 42168 38258 42180
rect 44910 42168 44916 42180
rect 44968 42168 44974 42220
rect 38838 42140 38844 42152
rect 35866 42112 38844 42140
rect 38838 42100 38844 42112
rect 38896 42100 38902 42152
rect 57422 41964 57428 42016
rect 57480 42004 57486 42016
rect 57885 42007 57943 42013
rect 57885 42004 57897 42007
rect 57480 41976 57897 42004
rect 57480 41964 57486 41976
rect 57885 41973 57897 41976
rect 57931 41973 57943 42007
rect 57885 41967 57943 41973
rect 1104 41914 68816 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 68816 41914
rect 1104 41840 68816 41862
rect 57422 41664 57428 41676
rect 57383 41636 57428 41664
rect 57422 41624 57428 41636
rect 57480 41624 57486 41676
rect 59078 41664 59084 41676
rect 59039 41636 59084 41664
rect 59078 41624 59084 41636
rect 59136 41624 59142 41676
rect 56778 41596 56784 41608
rect 56739 41568 56784 41596
rect 56778 41556 56784 41568
rect 56836 41556 56842 41608
rect 56873 41531 56931 41537
rect 56873 41497 56885 41531
rect 56919 41528 56931 41531
rect 57609 41531 57667 41537
rect 57609 41528 57621 41531
rect 56919 41500 57621 41528
rect 56919 41497 56931 41500
rect 56873 41491 56931 41497
rect 57609 41497 57621 41500
rect 57655 41497 57667 41531
rect 57609 41491 57667 41497
rect 1104 41370 68816 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 68816 41370
rect 1104 41296 68816 41318
rect 1104 40826 68816 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 68816 40826
rect 1104 40752 68816 40774
rect 1104 40282 68816 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 68816 40282
rect 1104 40208 68816 40230
rect 61378 40060 61384 40112
rect 61436 40100 61442 40112
rect 66162 40100 66168 40112
rect 61436 40072 66168 40100
rect 61436 40060 61442 40072
rect 66162 40060 66168 40072
rect 66220 40060 66226 40112
rect 9766 39788 9772 39840
rect 9824 39828 9830 39840
rect 9861 39831 9919 39837
rect 9861 39828 9873 39831
rect 9824 39800 9873 39828
rect 9824 39788 9830 39800
rect 9861 39797 9873 39800
rect 9907 39797 9919 39831
rect 9861 39791 9919 39797
rect 1104 39738 68816 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 68816 39738
rect 1104 39664 68816 39686
rect 6886 39528 10272 39556
rect 3602 39312 3608 39364
rect 3660 39352 3666 39364
rect 6886 39352 6914 39528
rect 9766 39488 9772 39500
rect 9727 39460 9772 39488
rect 9766 39448 9772 39460
rect 9824 39448 9830 39500
rect 10244 39497 10272 39528
rect 10229 39491 10287 39497
rect 10229 39457 10241 39491
rect 10275 39457 10287 39491
rect 10229 39451 10287 39457
rect 32950 39380 32956 39432
rect 33008 39420 33014 39432
rect 33045 39423 33103 39429
rect 33045 39420 33057 39423
rect 33008 39392 33057 39420
rect 33008 39380 33014 39392
rect 33045 39389 33057 39392
rect 33091 39389 33103 39423
rect 33045 39383 33103 39389
rect 3660 39324 6914 39352
rect 9953 39355 10011 39361
rect 3660 39312 3666 39324
rect 9953 39321 9965 39355
rect 9999 39352 10011 39355
rect 10410 39352 10416 39364
rect 9999 39324 10416 39352
rect 9999 39321 10011 39324
rect 9953 39315 10011 39321
rect 10410 39312 10416 39324
rect 10468 39312 10474 39364
rect 1104 39194 68816 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 68816 39194
rect 1104 39120 68816 39142
rect 10410 39080 10416 39092
rect 10371 39052 10416 39080
rect 10410 39040 10416 39052
rect 10468 39040 10474 39092
rect 64785 39015 64843 39021
rect 64785 38981 64797 39015
rect 64831 39012 64843 39015
rect 65521 39015 65579 39021
rect 65521 39012 65533 39015
rect 64831 38984 65533 39012
rect 64831 38981 64843 38984
rect 64785 38975 64843 38981
rect 65521 38981 65533 38984
rect 65567 38981 65579 39015
rect 65521 38975 65579 38981
rect 10502 38944 10508 38956
rect 10463 38916 10508 38944
rect 10502 38904 10508 38916
rect 10560 38904 10566 38956
rect 32950 38944 32956 38956
rect 32911 38916 32956 38944
rect 32950 38904 32956 38916
rect 33008 38904 33014 38956
rect 64690 38944 64696 38956
rect 64651 38916 64696 38944
rect 64690 38904 64696 38916
rect 64748 38904 64754 38956
rect 33134 38876 33140 38888
rect 33095 38848 33140 38876
rect 33134 38836 33140 38848
rect 33192 38836 33198 38888
rect 34793 38879 34851 38885
rect 34793 38845 34805 38879
rect 34839 38876 34851 38879
rect 65150 38876 65156 38888
rect 34839 38848 65156 38876
rect 34839 38845 34851 38848
rect 34793 38839 34851 38845
rect 65150 38836 65156 38848
rect 65208 38836 65214 38888
rect 65334 38876 65340 38888
rect 65295 38848 65340 38876
rect 65334 38836 65340 38848
rect 65392 38836 65398 38888
rect 67174 38876 67180 38888
rect 67135 38848 67180 38876
rect 67174 38836 67180 38848
rect 67232 38836 67238 38888
rect 1104 38650 68816 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 68816 38650
rect 1104 38576 68816 38598
rect 32953 38539 33011 38545
rect 32953 38505 32965 38539
rect 32999 38536 33011 38539
rect 33134 38536 33140 38548
rect 32999 38508 33140 38536
rect 32999 38505 33011 38508
rect 32953 38499 33011 38505
rect 33134 38496 33140 38508
rect 33192 38496 33198 38548
rect 65334 38496 65340 38548
rect 65392 38536 65398 38548
rect 65613 38539 65671 38545
rect 65613 38536 65625 38539
rect 65392 38508 65625 38536
rect 65392 38496 65398 38508
rect 65613 38505 65625 38508
rect 65659 38505 65671 38539
rect 65613 38499 65671 38505
rect 32858 38332 32864 38344
rect 32819 38304 32864 38332
rect 32858 38292 32864 38304
rect 32916 38292 32922 38344
rect 1104 38106 68816 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 68816 38106
rect 1104 38032 68816 38054
rect 37366 37652 37372 37664
rect 37327 37624 37372 37652
rect 37366 37612 37372 37624
rect 37424 37612 37430 37664
rect 61654 37652 61660 37664
rect 61615 37624 61660 37652
rect 61654 37612 61660 37624
rect 61712 37612 61718 37664
rect 1104 37562 68816 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 68816 37562
rect 1104 37488 68816 37510
rect 37366 37312 37372 37324
rect 37327 37284 37372 37312
rect 37366 37272 37372 37284
rect 37424 37272 37430 37324
rect 61654 37312 61660 37324
rect 61615 37284 61660 37312
rect 61654 37272 61660 37284
rect 61712 37272 61718 37324
rect 63497 37315 63555 37321
rect 63497 37281 63509 37315
rect 63543 37312 63555 37315
rect 66162 37312 66168 37324
rect 63543 37284 66168 37312
rect 63543 37281 63555 37284
rect 63497 37275 63555 37281
rect 66162 37272 66168 37284
rect 66220 37272 66226 37324
rect 35345 37247 35403 37253
rect 35345 37244 35357 37247
rect 32416 37216 35357 37244
rect 32416 37188 32444 37216
rect 35345 37213 35357 37216
rect 35391 37213 35403 37247
rect 39206 37244 39212 37256
rect 39167 37216 39212 37244
rect 35345 37207 35403 37213
rect 32398 37176 32404 37188
rect 32359 37148 32404 37176
rect 32398 37136 32404 37148
rect 32456 37136 32462 37188
rect 35360 37176 35388 37207
rect 39206 37204 39212 37216
rect 39264 37204 39270 37256
rect 60918 37204 60924 37256
rect 60976 37244 60982 37256
rect 61013 37247 61071 37253
rect 61013 37244 61025 37247
rect 60976 37216 61025 37244
rect 60976 37204 60982 37216
rect 61013 37213 61025 37216
rect 61059 37244 61071 37247
rect 61286 37244 61292 37256
rect 61059 37216 61292 37244
rect 61059 37213 61071 37216
rect 61013 37207 61071 37213
rect 61286 37204 61292 37216
rect 61344 37204 61350 37256
rect 36538 37176 36544 37188
rect 35360 37148 36544 37176
rect 36538 37136 36544 37148
rect 36596 37136 36602 37188
rect 36630 37136 36636 37188
rect 36688 37176 36694 37188
rect 37553 37179 37611 37185
rect 37553 37176 37565 37179
rect 36688 37148 37565 37176
rect 36688 37136 36694 37148
rect 37553 37145 37565 37148
rect 37599 37145 37611 37179
rect 37553 37139 37611 37145
rect 61105 37179 61163 37185
rect 61105 37145 61117 37179
rect 61151 37176 61163 37179
rect 61841 37179 61899 37185
rect 61841 37176 61853 37179
rect 61151 37148 61853 37176
rect 61151 37145 61163 37148
rect 61105 37139 61163 37145
rect 61841 37145 61853 37148
rect 61887 37145 61899 37179
rect 61841 37139 61899 37145
rect 32490 37108 32496 37120
rect 32451 37080 32496 37108
rect 32490 37068 32496 37080
rect 32548 37068 32554 37120
rect 35529 37111 35587 37117
rect 35529 37077 35541 37111
rect 35575 37108 35587 37111
rect 37366 37108 37372 37120
rect 35575 37080 37372 37108
rect 35575 37077 35587 37080
rect 35529 37071 35587 37077
rect 37366 37068 37372 37080
rect 37424 37068 37430 37120
rect 1104 37018 68816 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 68816 37018
rect 1104 36944 68816 36966
rect 36630 36904 36636 36916
rect 36591 36876 36636 36904
rect 36630 36864 36636 36876
rect 36688 36864 36694 36916
rect 38948 36876 45554 36904
rect 1578 36796 1584 36848
rect 1636 36836 1642 36848
rect 32398 36836 32404 36848
rect 1636 36808 32404 36836
rect 1636 36796 1642 36808
rect 32398 36796 32404 36808
rect 32456 36796 32462 36848
rect 32490 36796 32496 36848
rect 32548 36836 32554 36848
rect 35437 36839 35495 36845
rect 32548 36808 34100 36836
rect 32548 36796 32554 36808
rect 32416 36768 32444 36796
rect 34072 36777 34100 36808
rect 35437 36805 35449 36839
rect 35483 36836 35495 36839
rect 35618 36836 35624 36848
rect 35483 36808 35624 36836
rect 35483 36805 35495 36808
rect 35437 36799 35495 36805
rect 35618 36796 35624 36808
rect 35676 36796 35682 36848
rect 35728 36808 36584 36836
rect 33137 36771 33195 36777
rect 33137 36768 33149 36771
rect 32416 36740 33149 36768
rect 33137 36737 33149 36740
rect 33183 36737 33195 36771
rect 33137 36731 33195 36737
rect 34057 36771 34115 36777
rect 34057 36737 34069 36771
rect 34103 36737 34115 36771
rect 34057 36731 34115 36737
rect 34146 36728 34152 36780
rect 34204 36768 34210 36780
rect 35728 36768 35756 36808
rect 34204 36740 35756 36768
rect 35805 36771 35863 36777
rect 34204 36728 34210 36740
rect 35805 36737 35817 36771
rect 35851 36768 35863 36771
rect 36078 36768 36084 36780
rect 35851 36740 36084 36768
rect 35851 36737 35863 36740
rect 35805 36731 35863 36737
rect 36078 36728 36084 36740
rect 36136 36728 36142 36780
rect 36556 36777 36584 36808
rect 37642 36796 37648 36848
rect 37700 36836 37706 36848
rect 37918 36836 37924 36848
rect 37700 36808 37924 36836
rect 37700 36796 37706 36808
rect 37918 36796 37924 36808
rect 37976 36796 37982 36848
rect 38010 36796 38016 36848
rect 38068 36836 38074 36848
rect 38948 36845 38976 36876
rect 38933 36839 38991 36845
rect 38933 36836 38945 36839
rect 38068 36808 38945 36836
rect 38068 36796 38074 36808
rect 38933 36805 38945 36808
rect 38979 36805 38991 36839
rect 40310 36836 40316 36848
rect 40271 36808 40316 36836
rect 38933 36799 38991 36805
rect 40310 36796 40316 36808
rect 40368 36796 40374 36848
rect 36541 36771 36599 36777
rect 36541 36737 36553 36771
rect 36587 36737 36599 36771
rect 37366 36768 37372 36780
rect 37327 36740 37372 36768
rect 36541 36731 36599 36737
rect 37366 36728 37372 36740
rect 37424 36768 37430 36780
rect 38565 36771 38623 36777
rect 38565 36768 38577 36771
rect 37424 36740 38577 36768
rect 37424 36728 37430 36740
rect 38565 36737 38577 36740
rect 38611 36737 38623 36771
rect 38565 36731 38623 36737
rect 38654 36728 38660 36780
rect 38712 36768 38718 36780
rect 39761 36771 39819 36777
rect 39761 36768 39773 36771
rect 38712 36740 39773 36768
rect 38712 36728 38718 36740
rect 39761 36737 39773 36740
rect 39807 36737 39819 36771
rect 45526 36768 45554 36876
rect 64690 36768 64696 36780
rect 45526 36740 64696 36768
rect 39761 36731 39819 36737
rect 64690 36728 64696 36740
rect 64748 36768 64754 36780
rect 64785 36771 64843 36777
rect 64785 36768 64797 36771
rect 64748 36740 64797 36768
rect 64748 36728 64754 36740
rect 64785 36737 64797 36740
rect 64831 36737 64843 36771
rect 64785 36731 64843 36737
rect 13449 36703 13507 36709
rect 13449 36669 13461 36703
rect 13495 36700 13507 36703
rect 13909 36703 13967 36709
rect 13909 36700 13921 36703
rect 13495 36672 13921 36700
rect 13495 36669 13507 36672
rect 13449 36663 13507 36669
rect 13909 36669 13921 36672
rect 13955 36669 13967 36703
rect 13909 36663 13967 36669
rect 14093 36703 14151 36709
rect 14093 36669 14105 36703
rect 14139 36700 14151 36703
rect 14182 36700 14188 36712
rect 14139 36672 14188 36700
rect 14139 36669 14151 36672
rect 14093 36663 14151 36669
rect 14182 36660 14188 36672
rect 14240 36660 14246 36712
rect 14369 36703 14427 36709
rect 14369 36669 14381 36703
rect 14415 36669 14427 36703
rect 14369 36663 14427 36669
rect 34425 36703 34483 36709
rect 34425 36669 34437 36703
rect 34471 36700 34483 36703
rect 34698 36700 34704 36712
rect 34471 36672 34704 36700
rect 34471 36669 34483 36672
rect 34425 36663 34483 36669
rect 13814 36592 13820 36644
rect 13872 36632 13878 36644
rect 14384 36632 14412 36663
rect 34698 36660 34704 36672
rect 34756 36700 34762 36712
rect 35434 36700 35440 36712
rect 34756 36672 35440 36700
rect 34756 36660 34762 36672
rect 35434 36660 35440 36672
rect 35492 36660 35498 36712
rect 13872 36604 14412 36632
rect 13872 36592 13878 36604
rect 33413 36567 33471 36573
rect 33413 36533 33425 36567
rect 33459 36564 33471 36567
rect 34422 36564 34428 36576
rect 33459 36536 34428 36564
rect 33459 36533 33471 36536
rect 33413 36527 33471 36533
rect 34422 36524 34428 36536
rect 34480 36524 34486 36576
rect 64874 36524 64880 36576
rect 64932 36564 64938 36576
rect 64932 36536 64977 36564
rect 64932 36524 64938 36536
rect 65518 36524 65524 36576
rect 65576 36564 65582 36576
rect 65613 36567 65671 36573
rect 65613 36564 65625 36567
rect 65576 36536 65625 36564
rect 65576 36524 65582 36536
rect 65613 36533 65625 36536
rect 65659 36533 65671 36567
rect 65613 36527 65671 36533
rect 1104 36474 68816 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 68816 36474
rect 1104 36400 68816 36422
rect 14182 36360 14188 36372
rect 14143 36332 14188 36360
rect 14182 36320 14188 36332
rect 14240 36320 14246 36372
rect 32950 36320 32956 36372
rect 33008 36360 33014 36372
rect 43346 36360 43352 36372
rect 33008 36332 43352 36360
rect 33008 36320 33014 36332
rect 43346 36320 43352 36332
rect 43404 36320 43410 36372
rect 25314 36252 25320 36304
rect 25372 36292 25378 36304
rect 25372 36264 26234 36292
rect 25372 36252 25378 36264
rect 26206 36224 26234 36264
rect 64874 36252 64880 36304
rect 64932 36292 64938 36304
rect 64932 36264 65840 36292
rect 64932 36252 64938 36264
rect 38105 36227 38163 36233
rect 38105 36224 38117 36227
rect 26206 36196 38117 36224
rect 38105 36193 38117 36196
rect 38151 36224 38163 36227
rect 43438 36224 43444 36236
rect 38151 36196 43444 36224
rect 38151 36193 38163 36196
rect 38105 36187 38163 36193
rect 43438 36184 43444 36196
rect 43496 36184 43502 36236
rect 65518 36184 65524 36236
rect 65576 36224 65582 36236
rect 65812 36233 65840 36264
rect 65613 36227 65671 36233
rect 65613 36224 65625 36227
rect 65576 36196 65625 36224
rect 65576 36184 65582 36196
rect 65613 36193 65625 36196
rect 65659 36193 65671 36227
rect 65613 36187 65671 36193
rect 65797 36227 65855 36233
rect 65797 36193 65809 36227
rect 65843 36193 65855 36227
rect 65797 36187 65855 36193
rect 6362 36156 6368 36168
rect 6323 36128 6368 36156
rect 6362 36116 6368 36128
rect 6420 36116 6426 36168
rect 14274 36156 14280 36168
rect 14235 36128 14280 36156
rect 14274 36116 14280 36128
rect 14332 36116 14338 36168
rect 32401 36159 32459 36165
rect 32401 36125 32413 36159
rect 32447 36156 32459 36159
rect 32490 36156 32496 36168
rect 32447 36128 32496 36156
rect 32447 36125 32459 36128
rect 32401 36119 32459 36125
rect 32490 36116 32496 36128
rect 32548 36156 32554 36168
rect 33505 36159 33563 36165
rect 33505 36156 33517 36159
rect 32548 36128 33517 36156
rect 32548 36116 32554 36128
rect 33505 36125 33517 36128
rect 33551 36125 33563 36159
rect 33778 36156 33784 36168
rect 33691 36128 33784 36156
rect 33505 36119 33563 36125
rect 33778 36116 33784 36128
rect 33836 36156 33842 36168
rect 34146 36156 34152 36168
rect 33836 36128 34152 36156
rect 33836 36116 33842 36128
rect 34146 36116 34152 36128
rect 34204 36116 34210 36168
rect 36078 36156 36084 36168
rect 35991 36128 36084 36156
rect 36078 36116 36084 36128
rect 36136 36116 36142 36168
rect 36538 36156 36544 36168
rect 36499 36128 36544 36156
rect 36538 36116 36544 36128
rect 36596 36116 36602 36168
rect 37366 36116 37372 36168
rect 37424 36156 37430 36168
rect 37553 36159 37611 36165
rect 37553 36156 37565 36159
rect 37424 36128 37565 36156
rect 37424 36116 37430 36128
rect 37553 36125 37565 36128
rect 37599 36125 37611 36159
rect 37553 36119 37611 36125
rect 45186 36116 45192 36168
rect 45244 36156 45250 36168
rect 45373 36159 45431 36165
rect 45373 36156 45385 36159
rect 45244 36128 45385 36156
rect 45244 36116 45250 36128
rect 45373 36125 45385 36128
rect 45419 36125 45431 36159
rect 45373 36119 45431 36125
rect 32766 36048 32772 36100
rect 32824 36088 32830 36100
rect 32950 36088 32956 36100
rect 32824 36060 32956 36088
rect 32824 36048 32830 36060
rect 32950 36048 32956 36060
rect 33008 36048 33014 36100
rect 35253 36091 35311 36097
rect 35253 36057 35265 36091
rect 35299 36088 35311 36091
rect 35299 36060 35333 36088
rect 35299 36057 35311 36060
rect 35253 36051 35311 36057
rect 26234 35980 26240 36032
rect 26292 36020 26298 36032
rect 35268 36020 35296 36051
rect 35434 36020 35440 36032
rect 26292 35992 35440 36020
rect 26292 35980 26298 35992
rect 35434 35980 35440 35992
rect 35492 35980 35498 36032
rect 35894 35980 35900 36032
rect 35952 36020 35958 36032
rect 36096 36020 36124 36116
rect 67450 36088 67456 36100
rect 67411 36060 67456 36088
rect 67450 36048 67456 36060
rect 67508 36048 67514 36100
rect 36725 36023 36783 36029
rect 36725 36020 36737 36023
rect 35952 35992 36737 36020
rect 35952 35980 35958 35992
rect 36725 35989 36737 35992
rect 36771 35989 36783 36023
rect 36725 35983 36783 35989
rect 1104 35930 68816 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 68816 35930
rect 1104 35856 68816 35878
rect 34517 35751 34575 35757
rect 34517 35717 34529 35751
rect 34563 35748 34575 35751
rect 40678 35748 40684 35760
rect 34563 35720 40684 35748
rect 34563 35717 34575 35720
rect 34517 35711 34575 35717
rect 40678 35708 40684 35720
rect 40736 35708 40742 35760
rect 47029 35751 47087 35757
rect 47029 35717 47041 35751
rect 47075 35748 47087 35751
rect 61378 35748 61384 35760
rect 47075 35720 61384 35748
rect 47075 35717 47087 35720
rect 47029 35711 47087 35717
rect 61378 35708 61384 35720
rect 61436 35708 61442 35760
rect 6362 35680 6368 35692
rect 6323 35652 6368 35680
rect 6362 35640 6368 35652
rect 6420 35640 6426 35692
rect 32490 35640 32496 35692
rect 32548 35680 32554 35692
rect 32861 35683 32919 35689
rect 32861 35680 32873 35683
rect 32548 35652 32873 35680
rect 32548 35640 32554 35652
rect 32861 35649 32873 35652
rect 32907 35680 32919 35683
rect 33965 35683 34023 35689
rect 33965 35680 33977 35683
rect 32907 35652 33977 35680
rect 32907 35649 32919 35652
rect 32861 35643 32919 35649
rect 33965 35649 33977 35652
rect 34011 35649 34023 35683
rect 33965 35643 34023 35649
rect 35894 35640 35900 35692
rect 35952 35680 35958 35692
rect 35952 35652 35997 35680
rect 35952 35640 35958 35652
rect 41414 35640 41420 35692
rect 41472 35680 41478 35692
rect 44545 35683 44603 35689
rect 44545 35680 44557 35683
rect 41472 35652 44557 35680
rect 41472 35640 41478 35652
rect 44545 35649 44557 35652
rect 44591 35649 44603 35683
rect 45186 35680 45192 35692
rect 45147 35652 45192 35680
rect 44545 35643 44603 35649
rect 45186 35640 45192 35652
rect 45244 35640 45250 35692
rect 6546 35612 6552 35624
rect 6507 35584 6552 35612
rect 6546 35572 6552 35584
rect 6604 35572 6610 35624
rect 6825 35615 6883 35621
rect 6825 35581 6837 35615
rect 6871 35581 6883 35615
rect 6825 35575 6883 35581
rect 4062 35504 4068 35556
rect 4120 35544 4126 35556
rect 6840 35544 6868 35575
rect 14274 35572 14280 35624
rect 14332 35612 14338 35624
rect 32585 35615 32643 35621
rect 32585 35612 32597 35615
rect 14332 35584 32597 35612
rect 14332 35572 14338 35584
rect 32585 35581 32597 35584
rect 32631 35612 32643 35615
rect 34606 35612 34612 35624
rect 32631 35584 34612 35612
rect 32631 35581 32643 35584
rect 32585 35575 32643 35581
rect 34606 35572 34612 35584
rect 34664 35572 34670 35624
rect 35342 35612 35348 35624
rect 35303 35584 35348 35612
rect 35342 35572 35348 35584
rect 35400 35612 35406 35624
rect 44637 35615 44695 35621
rect 35400 35584 35894 35612
rect 35400 35572 35406 35584
rect 4120 35516 6868 35544
rect 35866 35544 35894 35584
rect 44637 35581 44649 35615
rect 44683 35612 44695 35615
rect 45373 35615 45431 35621
rect 45373 35612 45385 35615
rect 44683 35584 45385 35612
rect 44683 35581 44695 35584
rect 44637 35575 44695 35581
rect 45373 35581 45385 35584
rect 45419 35581 45431 35615
rect 61286 35612 61292 35624
rect 45373 35575 45431 35581
rect 55186 35584 61292 35612
rect 55186 35544 55214 35584
rect 61286 35572 61292 35584
rect 61344 35572 61350 35624
rect 35866 35516 55214 35544
rect 4120 35504 4126 35516
rect 1104 35386 68816 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 68816 35386
rect 1104 35312 68816 35334
rect 6457 35275 6515 35281
rect 6457 35241 6469 35275
rect 6503 35272 6515 35275
rect 6546 35272 6552 35284
rect 6503 35244 6552 35272
rect 6503 35241 6515 35244
rect 6457 35235 6515 35241
rect 6546 35232 6552 35244
rect 6604 35232 6610 35284
rect 6546 35068 6552 35080
rect 6507 35040 6552 35068
rect 6546 35028 6552 35040
rect 6604 35068 6610 35080
rect 14274 35068 14280 35080
rect 6604 35040 14280 35068
rect 6604 35028 6610 35040
rect 14274 35028 14280 35040
rect 14332 35028 14338 35080
rect 1104 34842 68816 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 68816 34842
rect 1104 34768 68816 34790
rect 34790 34552 34796 34604
rect 34848 34592 34854 34604
rect 35342 34592 35348 34604
rect 34848 34564 35348 34592
rect 34848 34552 34854 34564
rect 35342 34552 35348 34564
rect 35400 34552 35406 34604
rect 35894 34552 35900 34604
rect 35952 34592 35958 34604
rect 37366 34592 37372 34604
rect 35952 34564 35997 34592
rect 37327 34564 37372 34592
rect 35952 34552 35958 34564
rect 37366 34552 37372 34564
rect 37424 34552 37430 34604
rect 43254 34592 43260 34604
rect 37844 34564 43260 34592
rect 10502 34484 10508 34536
rect 10560 34524 10566 34536
rect 10962 34524 10968 34536
rect 10560 34496 10968 34524
rect 10560 34484 10566 34496
rect 10962 34484 10968 34496
rect 11020 34524 11026 34536
rect 35253 34527 35311 34533
rect 35253 34524 35265 34527
rect 11020 34496 35265 34524
rect 11020 34484 11026 34496
rect 35253 34493 35265 34496
rect 35299 34524 35311 34527
rect 37844 34524 37872 34564
rect 43254 34552 43260 34564
rect 43312 34552 43318 34604
rect 35299 34496 37872 34524
rect 37921 34527 37979 34533
rect 35299 34493 35311 34496
rect 35253 34487 35311 34493
rect 37921 34493 37933 34527
rect 37967 34524 37979 34527
rect 38194 34524 38200 34536
rect 37967 34496 38200 34524
rect 37967 34493 37979 34496
rect 37921 34487 37979 34493
rect 38194 34484 38200 34496
rect 38252 34484 38258 34536
rect 22002 34416 22008 34468
rect 22060 34456 22066 34468
rect 25314 34456 25320 34468
rect 22060 34428 25320 34456
rect 22060 34416 22066 34428
rect 25314 34416 25320 34428
rect 25372 34416 25378 34468
rect 24854 34388 24860 34400
rect 24815 34360 24860 34388
rect 24854 34348 24860 34360
rect 24912 34348 24918 34400
rect 1104 34298 68816 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 68816 34298
rect 1104 34224 68816 34246
rect 6886 34088 25360 34116
rect 3418 33872 3424 33924
rect 3476 33912 3482 33924
rect 6886 33912 6914 34088
rect 24854 34048 24860 34060
rect 24815 34020 24860 34048
rect 24854 34008 24860 34020
rect 24912 34008 24918 34060
rect 25332 34057 25360 34088
rect 25317 34051 25375 34057
rect 25317 34017 25329 34051
rect 25363 34017 25375 34051
rect 25317 34011 25375 34017
rect 35437 34051 35495 34057
rect 35437 34017 35449 34051
rect 35483 34048 35495 34051
rect 35526 34048 35532 34060
rect 35483 34020 35532 34048
rect 35483 34017 35495 34020
rect 35437 34011 35495 34017
rect 35526 34008 35532 34020
rect 35584 34008 35590 34060
rect 36446 34008 36452 34060
rect 36504 34048 36510 34060
rect 36725 34051 36783 34057
rect 36725 34048 36737 34051
rect 36504 34020 36737 34048
rect 36504 34008 36510 34020
rect 36725 34017 36737 34020
rect 36771 34048 36783 34051
rect 41414 34048 41420 34060
rect 36771 34020 41420 34048
rect 36771 34017 36783 34020
rect 36725 34011 36783 34017
rect 41414 34008 41420 34020
rect 41472 34008 41478 34060
rect 35713 33983 35771 33989
rect 35713 33949 35725 33983
rect 35759 33980 35771 33983
rect 35894 33980 35900 33992
rect 35759 33952 35900 33980
rect 35759 33949 35771 33952
rect 35713 33943 35771 33949
rect 35894 33940 35900 33952
rect 35952 33940 35958 33992
rect 37001 33983 37059 33989
rect 37001 33949 37013 33983
rect 37047 33980 37059 33983
rect 37366 33980 37372 33992
rect 37047 33952 37372 33980
rect 37047 33949 37059 33952
rect 37001 33943 37059 33949
rect 37366 33940 37372 33952
rect 37424 33940 37430 33992
rect 49142 33940 49148 33992
rect 49200 33980 49206 33992
rect 49237 33983 49295 33989
rect 49237 33980 49249 33983
rect 49200 33952 49249 33980
rect 49200 33940 49206 33952
rect 49237 33949 49249 33952
rect 49283 33949 49295 33983
rect 49237 33943 49295 33949
rect 55490 33940 55496 33992
rect 55548 33980 55554 33992
rect 55861 33983 55919 33989
rect 55861 33980 55873 33983
rect 55548 33952 55873 33980
rect 55548 33940 55554 33952
rect 55861 33949 55873 33952
rect 55907 33949 55919 33983
rect 55861 33943 55919 33949
rect 3476 33884 6914 33912
rect 25041 33915 25099 33921
rect 3476 33872 3482 33884
rect 25041 33881 25053 33915
rect 25087 33912 25099 33915
rect 25222 33912 25228 33924
rect 25087 33884 25228 33912
rect 25087 33881 25099 33884
rect 25041 33875 25099 33881
rect 25222 33872 25228 33884
rect 25280 33872 25286 33924
rect 1104 33754 68816 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 68816 33754
rect 1104 33680 68816 33702
rect 25222 33640 25228 33652
rect 25183 33612 25228 33640
rect 25222 33600 25228 33612
rect 25280 33600 25286 33652
rect 43346 33572 43352 33584
rect 41708 33544 43352 33572
rect 25314 33504 25320 33516
rect 25275 33476 25320 33504
rect 25314 33464 25320 33476
rect 25372 33464 25378 33516
rect 41708 33513 41736 33544
rect 43346 33532 43352 33544
rect 43404 33532 43410 33584
rect 66070 33572 66076 33584
rect 45526 33544 66076 33572
rect 41693 33507 41751 33513
rect 41693 33473 41705 33507
rect 41739 33473 41751 33507
rect 41693 33467 41751 33473
rect 42426 33436 42432 33448
rect 42387 33408 42432 33436
rect 42426 33396 42432 33408
rect 42484 33396 42490 33448
rect 42613 33439 42671 33445
rect 42613 33405 42625 33439
rect 42659 33405 42671 33439
rect 42613 33399 42671 33405
rect 44269 33439 44327 33445
rect 44269 33405 44281 33439
rect 44315 33436 44327 33439
rect 45526 33436 45554 33544
rect 66070 33532 66076 33544
rect 66128 33532 66134 33584
rect 49142 33504 49148 33516
rect 49103 33476 49148 33504
rect 49142 33464 49148 33476
rect 49200 33464 49206 33516
rect 55490 33504 55496 33516
rect 55451 33476 55496 33504
rect 55490 33464 55496 33476
rect 55548 33464 55554 33516
rect 49326 33436 49332 33448
rect 44315 33408 45554 33436
rect 49287 33408 49332 33436
rect 44315 33405 44327 33408
rect 44269 33399 44327 33405
rect 41785 33371 41843 33377
rect 41785 33337 41797 33371
rect 41831 33368 41843 33371
rect 42628 33368 42656 33399
rect 49326 33396 49332 33408
rect 49384 33396 49390 33448
rect 50985 33439 51043 33445
rect 50985 33405 50997 33439
rect 51031 33436 51043 33439
rect 55674 33436 55680 33448
rect 51031 33408 55214 33436
rect 55635 33408 55680 33436
rect 51031 33405 51043 33408
rect 50985 33399 51043 33405
rect 41831 33340 42656 33368
rect 55186 33368 55214 33408
rect 55674 33396 55680 33408
rect 55732 33396 55738 33448
rect 57330 33436 57336 33448
rect 57291 33408 57336 33436
rect 57330 33396 57336 33408
rect 57388 33396 57394 33448
rect 66162 33368 66168 33380
rect 55186 33340 66168 33368
rect 41831 33337 41843 33340
rect 41785 33331 41843 33337
rect 66162 33328 66168 33340
rect 66220 33328 66226 33380
rect 1104 33210 68816 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 68816 33210
rect 1104 33136 68816 33158
rect 42245 33099 42303 33105
rect 42245 33065 42257 33099
rect 42291 33096 42303 33099
rect 42426 33096 42432 33108
rect 42291 33068 42432 33096
rect 42291 33065 42303 33068
rect 42245 33059 42303 33065
rect 42426 33056 42432 33068
rect 42484 33056 42490 33108
rect 49145 33099 49203 33105
rect 49145 33065 49157 33099
rect 49191 33096 49203 33099
rect 49326 33096 49332 33108
rect 49191 33068 49332 33096
rect 49191 33065 49203 33068
rect 49145 33059 49203 33065
rect 49326 33056 49332 33068
rect 49384 33056 49390 33108
rect 55674 33056 55680 33108
rect 55732 33096 55738 33108
rect 56137 33099 56195 33105
rect 56137 33096 56149 33099
rect 55732 33068 56149 33096
rect 55732 33056 55738 33068
rect 56137 33065 56149 33068
rect 56183 33065 56195 33099
rect 56137 33059 56195 33065
rect 45526 32932 55214 32960
rect 40310 32852 40316 32904
rect 40368 32892 40374 32904
rect 45526 32892 45554 32932
rect 49050 32892 49056 32904
rect 40368 32864 45554 32892
rect 49011 32864 49056 32892
rect 40368 32852 40374 32864
rect 49050 32852 49056 32864
rect 49108 32852 49114 32904
rect 55186 32892 55214 32932
rect 56229 32895 56287 32901
rect 56229 32892 56241 32895
rect 55186 32864 56241 32892
rect 56229 32861 56241 32864
rect 56275 32861 56287 32895
rect 56229 32855 56287 32861
rect 1104 32666 68816 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 68816 32666
rect 1104 32592 68816 32614
rect 49050 32552 49056 32564
rect 43916 32524 49056 32552
rect 43438 32376 43444 32428
rect 43496 32416 43502 32428
rect 43916 32425 43944 32524
rect 49050 32512 49056 32524
rect 49108 32512 49114 32564
rect 43993 32487 44051 32493
rect 43993 32453 44005 32487
rect 44039 32484 44051 32487
rect 44729 32487 44787 32493
rect 44729 32484 44741 32487
rect 44039 32456 44741 32484
rect 44039 32453 44051 32456
rect 43993 32447 44051 32453
rect 44729 32453 44741 32456
rect 44775 32453 44787 32487
rect 44729 32447 44787 32453
rect 43901 32419 43959 32425
rect 43901 32416 43913 32419
rect 43496 32388 43913 32416
rect 43496 32376 43502 32388
rect 43901 32385 43913 32388
rect 43947 32385 43959 32419
rect 43901 32379 43959 32385
rect 44542 32348 44548 32360
rect 44503 32320 44548 32348
rect 44542 32308 44548 32320
rect 44600 32308 44606 32360
rect 45005 32351 45063 32357
rect 45005 32317 45017 32351
rect 45051 32317 45063 32351
rect 45005 32311 45063 32317
rect 44174 32240 44180 32292
rect 44232 32280 44238 32292
rect 45020 32280 45048 32311
rect 44232 32252 45048 32280
rect 44232 32240 44238 32252
rect 1104 32122 68816 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 68816 32122
rect 1104 32048 68816 32070
rect 44542 31968 44548 32020
rect 44600 32008 44606 32020
rect 45005 32011 45063 32017
rect 45005 32008 45017 32011
rect 44600 31980 45017 32008
rect 44600 31968 44606 31980
rect 45005 31977 45017 31980
rect 45051 31977 45063 32011
rect 45005 31971 45063 31977
rect 5442 31804 5448 31816
rect 5403 31776 5448 31804
rect 5442 31764 5448 31776
rect 5500 31764 5506 31816
rect 1104 31578 68816 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 68816 31578
rect 1104 31504 68816 31526
rect 6546 31328 6552 31340
rect 6507 31300 6552 31328
rect 6546 31288 6552 31300
rect 6604 31288 6610 31340
rect 34422 31288 34428 31340
rect 34480 31328 34486 31340
rect 38289 31331 38347 31337
rect 38289 31328 38301 31331
rect 34480 31300 38301 31328
rect 34480 31288 34486 31300
rect 38289 31297 38301 31300
rect 38335 31328 38347 31331
rect 38562 31328 38568 31340
rect 38335 31300 38568 31328
rect 38335 31297 38347 31300
rect 38289 31291 38347 31297
rect 38562 31288 38568 31300
rect 38620 31288 38626 31340
rect 38838 31260 38844 31272
rect 38799 31232 38844 31260
rect 38838 31220 38844 31232
rect 38896 31260 38902 31272
rect 56778 31260 56784 31272
rect 38896 31232 56784 31260
rect 38896 31220 38902 31232
rect 56778 31220 56784 31232
rect 56836 31260 56842 31272
rect 58158 31260 58164 31272
rect 56836 31232 58164 31260
rect 56836 31220 56842 31232
rect 58158 31220 58164 31232
rect 58216 31220 58222 31272
rect 5626 31084 5632 31136
rect 5684 31124 5690 31136
rect 6457 31127 6515 31133
rect 6457 31124 6469 31127
rect 5684 31096 6469 31124
rect 5684 31084 5690 31096
rect 6457 31093 6469 31096
rect 6503 31093 6515 31127
rect 6457 31087 6515 31093
rect 1104 31034 68816 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 68816 31034
rect 1104 30960 68816 30982
rect 2958 30812 2964 30864
rect 3016 30852 3022 30864
rect 3016 30824 5948 30852
rect 3016 30812 3022 30824
rect 5442 30784 5448 30796
rect 5403 30756 5448 30784
rect 5442 30744 5448 30756
rect 5500 30744 5506 30796
rect 5626 30784 5632 30796
rect 5587 30756 5632 30784
rect 5626 30744 5632 30756
rect 5684 30744 5690 30796
rect 5920 30793 5948 30824
rect 5905 30787 5963 30793
rect 5905 30753 5917 30787
rect 5951 30753 5963 30787
rect 32858 30784 32864 30796
rect 32819 30756 32864 30784
rect 5905 30747 5963 30753
rect 32858 30744 32864 30756
rect 32916 30744 32922 30796
rect 7742 30676 7748 30728
rect 7800 30716 7806 30728
rect 7837 30719 7895 30725
rect 7837 30716 7849 30719
rect 7800 30688 7849 30716
rect 7800 30676 7806 30688
rect 7837 30685 7849 30688
rect 7883 30685 7895 30719
rect 7837 30679 7895 30685
rect 19426 30676 19432 30728
rect 19484 30716 19490 30728
rect 19521 30719 19579 30725
rect 19521 30716 19533 30719
rect 19484 30688 19533 30716
rect 19484 30676 19490 30688
rect 19521 30685 19533 30688
rect 19567 30685 19579 30719
rect 19521 30679 19579 30685
rect 27982 30676 27988 30728
rect 28040 30716 28046 30728
rect 28077 30719 28135 30725
rect 28077 30716 28089 30719
rect 28040 30688 28089 30716
rect 28040 30676 28046 30688
rect 28077 30685 28089 30688
rect 28123 30685 28135 30719
rect 28077 30679 28135 30685
rect 33413 30719 33471 30725
rect 33413 30685 33425 30719
rect 33459 30716 33471 30719
rect 33594 30716 33600 30728
rect 33459 30688 33600 30716
rect 33459 30685 33471 30688
rect 33413 30679 33471 30685
rect 33594 30676 33600 30688
rect 33652 30716 33658 30728
rect 34422 30716 34428 30728
rect 33652 30688 34428 30716
rect 33652 30676 33658 30688
rect 34422 30676 34428 30688
rect 34480 30676 34486 30728
rect 59722 30716 59728 30728
rect 59683 30688 59728 30716
rect 59722 30676 59728 30688
rect 59780 30676 59786 30728
rect 60458 30716 60464 30728
rect 60419 30688 60464 30716
rect 60458 30676 60464 30688
rect 60516 30676 60522 30728
rect 59817 30651 59875 30657
rect 59817 30617 59829 30651
rect 59863 30648 59875 30651
rect 60645 30651 60703 30657
rect 60645 30648 60657 30651
rect 59863 30620 60657 30648
rect 59863 30617 59875 30620
rect 59817 30611 59875 30617
rect 60645 30617 60657 30620
rect 60691 30617 60703 30651
rect 60645 30611 60703 30617
rect 62301 30651 62359 30657
rect 62301 30617 62313 30651
rect 62347 30648 62359 30651
rect 66162 30648 66168 30660
rect 62347 30620 66168 30648
rect 62347 30617 62359 30620
rect 62301 30611 62359 30617
rect 66162 30608 66168 30620
rect 66220 30608 66226 30660
rect 1104 30490 68816 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 68816 30490
rect 1104 30416 68816 30438
rect 7742 30240 7748 30252
rect 7703 30212 7748 30240
rect 7742 30200 7748 30212
rect 7800 30200 7806 30252
rect 19426 30240 19432 30252
rect 19387 30212 19432 30240
rect 19426 30200 19432 30212
rect 19484 30200 19490 30252
rect 26145 30243 26203 30249
rect 26145 30209 26157 30243
rect 26191 30240 26203 30243
rect 27798 30240 27804 30252
rect 26191 30212 27804 30240
rect 26191 30209 26203 30212
rect 26145 30203 26203 30209
rect 27798 30200 27804 30212
rect 27856 30200 27862 30252
rect 27982 30240 27988 30252
rect 27943 30212 27988 30240
rect 27982 30200 27988 30212
rect 28040 30200 28046 30252
rect 60185 30243 60243 30249
rect 60185 30209 60197 30243
rect 60231 30240 60243 30243
rect 60458 30240 60464 30252
rect 60231 30212 60464 30240
rect 60231 30209 60243 30212
rect 60185 30203 60243 30209
rect 60458 30200 60464 30212
rect 60516 30200 60522 30252
rect 7929 30175 7987 30181
rect 7929 30141 7941 30175
rect 7975 30172 7987 30175
rect 8294 30172 8300 30184
rect 7975 30144 8300 30172
rect 7975 30141 7987 30144
rect 7929 30135 7987 30141
rect 8294 30132 8300 30144
rect 8352 30132 8358 30184
rect 8389 30175 8447 30181
rect 8389 30141 8401 30175
rect 8435 30141 8447 30175
rect 8389 30135 8447 30141
rect 19613 30175 19671 30181
rect 19613 30141 19625 30175
rect 19659 30172 19671 30175
rect 19978 30172 19984 30184
rect 19659 30144 19984 30172
rect 19659 30141 19671 30144
rect 19613 30135 19671 30141
rect 3602 30064 3608 30116
rect 3660 30104 3666 30116
rect 8404 30104 8432 30135
rect 19978 30132 19984 30144
rect 20036 30132 20042 30184
rect 20073 30175 20131 30181
rect 20073 30141 20085 30175
rect 20119 30141 20131 30175
rect 20073 30135 20131 30141
rect 28169 30175 28227 30181
rect 28169 30141 28181 30175
rect 28215 30172 28227 30175
rect 28350 30172 28356 30184
rect 28215 30144 28356 30172
rect 28215 30141 28227 30144
rect 28169 30135 28227 30141
rect 3660 30076 8432 30104
rect 3660 30064 3666 30076
rect 19334 30064 19340 30116
rect 19392 30104 19398 30116
rect 20088 30104 20116 30135
rect 28350 30132 28356 30144
rect 28408 30132 28414 30184
rect 28445 30175 28503 30181
rect 28445 30141 28457 30175
rect 28491 30141 28503 30175
rect 28445 30135 28503 30141
rect 19392 30076 20116 30104
rect 19392 30064 19398 30076
rect 26234 30064 26240 30116
rect 26292 30104 26298 30116
rect 28460 30104 28488 30135
rect 26292 30076 28488 30104
rect 26292 30064 26298 30076
rect 25498 30036 25504 30048
rect 25459 30008 25504 30036
rect 25498 29996 25504 30008
rect 25556 29996 25562 30048
rect 25682 29996 25688 30048
rect 25740 30036 25746 30048
rect 26053 30039 26111 30045
rect 26053 30036 26065 30039
rect 25740 30008 26065 30036
rect 25740 29996 25746 30008
rect 26053 30005 26065 30008
rect 26099 30005 26111 30039
rect 27522 30036 27528 30048
rect 27483 30008 27528 30036
rect 26053 29999 26111 30005
rect 27522 29996 27528 30008
rect 27580 29996 27586 30048
rect 51074 29996 51080 30048
rect 51132 30036 51138 30048
rect 51169 30039 51227 30045
rect 51169 30036 51181 30039
rect 51132 30008 51181 30036
rect 51132 29996 51138 30008
rect 51169 30005 51181 30008
rect 51215 30005 51227 30039
rect 51169 29999 51227 30005
rect 1104 29946 68816 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 68816 29946
rect 1104 29872 68816 29894
rect 8294 29832 8300 29844
rect 8255 29804 8300 29832
rect 8294 29792 8300 29804
rect 8352 29792 8358 29844
rect 19978 29832 19984 29844
rect 19939 29804 19984 29832
rect 19978 29792 19984 29804
rect 20036 29792 20042 29844
rect 23474 29792 23480 29844
rect 23532 29832 23538 29844
rect 28350 29832 28356 29844
rect 23532 29804 26004 29832
rect 28311 29804 28356 29832
rect 23532 29792 23538 29804
rect 25498 29696 25504 29708
rect 25459 29668 25504 29696
rect 25498 29656 25504 29668
rect 25556 29656 25562 29708
rect 25682 29696 25688 29708
rect 25643 29668 25688 29696
rect 25682 29656 25688 29668
rect 25740 29656 25746 29708
rect 25976 29705 26004 29804
rect 28350 29792 28356 29804
rect 28408 29792 28414 29844
rect 26050 29724 26056 29776
rect 26108 29764 26114 29776
rect 32766 29764 32772 29776
rect 26108 29736 32772 29764
rect 26108 29724 26114 29736
rect 32766 29724 32772 29736
rect 32824 29724 32830 29776
rect 25961 29699 26019 29705
rect 25961 29665 25973 29699
rect 26007 29665 26019 29699
rect 25961 29659 26019 29665
rect 27798 29656 27804 29708
rect 27856 29696 27862 29708
rect 37642 29696 37648 29708
rect 27856 29668 37648 29696
rect 27856 29656 27862 29668
rect 8386 29628 8392 29640
rect 8347 29600 8392 29628
rect 8386 29588 8392 29600
rect 8444 29588 8450 29640
rect 28460 29637 28488 29668
rect 37642 29656 37648 29668
rect 37700 29656 37706 29708
rect 20073 29631 20131 29637
rect 20073 29597 20085 29631
rect 20119 29597 20131 29631
rect 20073 29591 20131 29597
rect 28445 29631 28503 29637
rect 28445 29597 28457 29631
rect 28491 29597 28503 29631
rect 28445 29591 28503 29597
rect 20088 29560 20116 29591
rect 35618 29588 35624 29640
rect 35676 29628 35682 29640
rect 50893 29631 50951 29637
rect 50893 29628 50905 29631
rect 35676 29600 50905 29628
rect 35676 29588 35682 29600
rect 50893 29597 50905 29600
rect 50939 29597 50951 29631
rect 50893 29591 50951 29597
rect 50982 29588 50988 29640
rect 51040 29628 51046 29640
rect 51537 29631 51595 29637
rect 51537 29628 51549 29631
rect 51040 29600 51549 29628
rect 51040 29588 51046 29600
rect 51537 29597 51549 29600
rect 51583 29597 51595 29631
rect 51537 29591 51595 29597
rect 26050 29560 26056 29572
rect 20088 29532 26056 29560
rect 26050 29520 26056 29532
rect 26108 29520 26114 29572
rect 51718 29560 51724 29572
rect 51679 29532 51724 29560
rect 51718 29520 51724 29532
rect 51776 29520 51782 29572
rect 53374 29560 53380 29572
rect 53335 29532 53380 29560
rect 53374 29520 53380 29532
rect 53432 29520 53438 29572
rect 50985 29495 51043 29501
rect 50985 29461 50997 29495
rect 51031 29492 51043 29495
rect 51258 29492 51264 29504
rect 51031 29464 51264 29492
rect 51031 29461 51043 29464
rect 50985 29455 51043 29461
rect 51258 29452 51264 29464
rect 51316 29452 51322 29504
rect 1104 29402 68816 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 68816 29402
rect 1104 29328 68816 29350
rect 35434 29248 35440 29300
rect 35492 29288 35498 29300
rect 35492 29260 38608 29288
rect 35492 29248 35498 29260
rect 17954 29180 17960 29232
rect 18012 29220 18018 29232
rect 38580 29220 38608 29260
rect 38654 29248 38660 29300
rect 38712 29288 38718 29300
rect 59722 29288 59728 29300
rect 38712 29260 59728 29288
rect 38712 29248 38718 29260
rect 59722 29248 59728 29260
rect 59780 29248 59786 29300
rect 51537 29223 51595 29229
rect 18012 29192 26234 29220
rect 38580 29192 45554 29220
rect 18012 29180 18018 29192
rect 26206 29016 26234 29192
rect 27522 29152 27528 29164
rect 27483 29124 27528 29152
rect 27522 29112 27528 29124
rect 27580 29112 27586 29164
rect 33778 29112 33784 29164
rect 33836 29152 33842 29164
rect 37369 29155 37427 29161
rect 37369 29152 37381 29155
rect 33836 29124 37381 29152
rect 33836 29112 33842 29124
rect 37369 29121 37381 29124
rect 37415 29121 37427 29155
rect 37369 29115 37427 29121
rect 37660 29124 38056 29152
rect 27706 29084 27712 29096
rect 27667 29056 27712 29084
rect 27706 29044 27712 29056
rect 27764 29044 27770 29096
rect 27985 29087 28043 29093
rect 27985 29053 27997 29087
rect 28031 29053 28043 29087
rect 27985 29047 28043 29053
rect 28000 29016 28028 29047
rect 30742 29044 30748 29096
rect 30800 29084 30806 29096
rect 37660 29084 37688 29124
rect 30800 29056 37688 29084
rect 37829 29087 37887 29093
rect 30800 29044 30806 29056
rect 37829 29053 37841 29087
rect 37875 29053 37887 29087
rect 38028 29084 38056 29124
rect 38562 29112 38568 29164
rect 38620 29152 38626 29164
rect 39117 29155 39175 29161
rect 39117 29152 39129 29155
rect 38620 29124 39129 29152
rect 38620 29112 38626 29124
rect 39117 29121 39129 29124
rect 39163 29121 39175 29155
rect 45526 29152 45554 29192
rect 51537 29189 51549 29223
rect 51583 29220 51595 29223
rect 51718 29220 51724 29232
rect 51583 29192 51724 29220
rect 51583 29189 51595 29192
rect 51537 29183 51595 29189
rect 51718 29180 51724 29192
rect 51776 29180 51782 29232
rect 51445 29155 51503 29161
rect 51445 29152 51457 29155
rect 45526 29124 51457 29152
rect 39117 29115 39175 29121
rect 51445 29121 51457 29124
rect 51491 29121 51503 29155
rect 51445 29115 51503 29121
rect 38841 29087 38899 29093
rect 38841 29084 38853 29087
rect 38028 29056 38853 29084
rect 37829 29047 37887 29053
rect 38841 29053 38853 29056
rect 38887 29084 38899 29087
rect 61654 29084 61660 29096
rect 38887 29056 61660 29084
rect 38887 29053 38899 29056
rect 38841 29047 38899 29053
rect 26206 28988 28028 29016
rect 28074 28976 28080 29028
rect 28132 29016 28138 29028
rect 37844 29016 37872 29047
rect 61654 29044 61660 29056
rect 61712 29044 61718 29096
rect 38654 29016 38660 29028
rect 28132 28988 38660 29016
rect 28132 28976 28138 28988
rect 38654 28976 38660 28988
rect 38712 28976 38718 29028
rect 50982 29016 50988 29028
rect 50943 28988 50988 29016
rect 50982 28976 50988 28988
rect 51040 28976 51046 29028
rect 3418 28908 3424 28960
rect 3476 28948 3482 28960
rect 23474 28948 23480 28960
rect 3476 28920 23480 28948
rect 3476 28908 3482 28920
rect 23474 28908 23480 28920
rect 23532 28908 23538 28960
rect 1104 28858 68816 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 68816 28858
rect 1104 28784 68816 28806
rect 27706 28704 27712 28756
rect 27764 28744 27770 28756
rect 28077 28747 28135 28753
rect 28077 28744 28089 28747
rect 27764 28716 28089 28744
rect 27764 28704 27770 28716
rect 28077 28713 28089 28716
rect 28123 28713 28135 28747
rect 28077 28707 28135 28713
rect 51074 28608 51080 28620
rect 51035 28580 51080 28608
rect 51074 28568 51080 28580
rect 51132 28568 51138 28620
rect 51258 28608 51264 28620
rect 51219 28580 51264 28608
rect 51258 28568 51264 28580
rect 51316 28568 51322 28620
rect 28169 28543 28227 28549
rect 28169 28509 28181 28543
rect 28215 28540 28227 28543
rect 30742 28540 30748 28552
rect 28215 28512 30748 28540
rect 28215 28509 28227 28512
rect 28169 28503 28227 28509
rect 30742 28500 30748 28512
rect 30800 28500 30806 28552
rect 33594 28540 33600 28552
rect 33555 28512 33600 28540
rect 33594 28500 33600 28512
rect 33652 28500 33658 28552
rect 60642 28500 60648 28552
rect 60700 28540 60706 28552
rect 61197 28543 61255 28549
rect 61197 28540 61209 28543
rect 60700 28512 61209 28540
rect 60700 28500 60706 28512
rect 61197 28509 61209 28512
rect 61243 28509 61255 28543
rect 61197 28503 61255 28509
rect 8386 28432 8392 28484
rect 8444 28472 8450 28484
rect 9122 28472 9128 28484
rect 8444 28444 9128 28472
rect 8444 28432 8450 28444
rect 9122 28432 9128 28444
rect 9180 28472 9186 28484
rect 33137 28475 33195 28481
rect 33137 28472 33149 28475
rect 9180 28444 33149 28472
rect 9180 28432 9186 28444
rect 33137 28441 33149 28444
rect 33183 28472 33195 28475
rect 40126 28472 40132 28484
rect 33183 28444 40132 28472
rect 33183 28441 33195 28444
rect 33137 28435 33195 28441
rect 40126 28432 40132 28444
rect 40184 28432 40190 28484
rect 52914 28472 52920 28484
rect 52875 28444 52920 28472
rect 52914 28432 52920 28444
rect 52972 28432 52978 28484
rect 1104 28314 68816 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 68816 28314
rect 1104 28240 68816 28262
rect 60642 28064 60648 28076
rect 60603 28036 60648 28064
rect 60642 28024 60648 28036
rect 60700 28024 60706 28076
rect 49881 27999 49939 28005
rect 49881 27965 49893 27999
rect 49927 27996 49939 27999
rect 50341 27999 50399 28005
rect 50341 27996 50353 27999
rect 49927 27968 50353 27996
rect 49927 27965 49939 27968
rect 49881 27959 49939 27965
rect 50341 27965 50353 27968
rect 50387 27965 50399 27999
rect 50522 27996 50528 28008
rect 50483 27968 50528 27996
rect 50341 27959 50399 27965
rect 50522 27956 50528 27968
rect 50580 27956 50586 28008
rect 52181 27999 52239 28005
rect 52181 27965 52193 27999
rect 52227 27996 52239 27999
rect 60826 27996 60832 28008
rect 52227 27968 55214 27996
rect 60787 27968 60832 27996
rect 52227 27965 52239 27968
rect 52181 27959 52239 27965
rect 55186 27928 55214 27968
rect 60826 27956 60832 27968
rect 60884 27956 60890 28008
rect 62485 27999 62543 28005
rect 62485 27965 62497 27999
rect 62531 27996 62543 27999
rect 64966 27996 64972 28008
rect 62531 27968 64972 27996
rect 62531 27965 62543 27968
rect 62485 27959 62543 27965
rect 64966 27956 64972 27968
rect 65024 27956 65030 28008
rect 66162 27928 66168 27940
rect 55186 27900 66168 27928
rect 66162 27888 66168 27900
rect 66220 27888 66226 27940
rect 1104 27770 68816 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 68816 27770
rect 1104 27696 68816 27718
rect 50522 27656 50528 27668
rect 50483 27628 50528 27656
rect 50522 27616 50528 27628
rect 50580 27616 50586 27668
rect 60826 27616 60832 27668
rect 60884 27656 60890 27668
rect 61197 27659 61255 27665
rect 61197 27656 61209 27659
rect 60884 27628 61209 27656
rect 60884 27616 60890 27628
rect 61197 27625 61209 27628
rect 61243 27625 61255 27659
rect 61197 27619 61255 27625
rect 34698 27548 34704 27600
rect 34756 27588 34762 27600
rect 35342 27588 35348 27600
rect 34756 27560 35348 27588
rect 34756 27548 34762 27560
rect 35342 27548 35348 27560
rect 35400 27548 35406 27600
rect 35526 27412 35532 27464
rect 35584 27452 35590 27464
rect 50433 27455 50491 27461
rect 50433 27452 50445 27455
rect 35584 27424 50445 27452
rect 35584 27412 35590 27424
rect 50433 27421 50445 27424
rect 50479 27421 50491 27455
rect 61286 27452 61292 27464
rect 61247 27424 61292 27452
rect 50433 27415 50491 27421
rect 61286 27412 61292 27424
rect 61344 27412 61350 27464
rect 1104 27226 68816 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 68816 27226
rect 1104 27152 68816 27174
rect 33778 26908 33784 26920
rect 33739 26880 33784 26908
rect 33778 26868 33784 26880
rect 33836 26868 33842 26920
rect 33965 26911 34023 26917
rect 33965 26877 33977 26911
rect 34011 26908 34023 26911
rect 34790 26908 34796 26920
rect 34011 26880 34796 26908
rect 34011 26877 34023 26880
rect 33965 26871 34023 26877
rect 34790 26868 34796 26880
rect 34848 26868 34854 26920
rect 34885 26911 34943 26917
rect 34885 26877 34897 26911
rect 34931 26877 34943 26911
rect 34885 26871 34943 26877
rect 6914 26800 6920 26852
rect 6972 26840 6978 26852
rect 34900 26840 34928 26871
rect 6972 26812 34928 26840
rect 6972 26800 6978 26812
rect 55766 26732 55772 26784
rect 55824 26772 55830 26784
rect 56413 26775 56471 26781
rect 56413 26772 56425 26775
rect 55824 26744 56425 26772
rect 55824 26732 55830 26744
rect 56413 26741 56425 26744
rect 56459 26741 56471 26775
rect 56413 26735 56471 26741
rect 58066 26732 58072 26784
rect 58124 26772 58130 26784
rect 58253 26775 58311 26781
rect 58253 26772 58265 26775
rect 58124 26744 58265 26772
rect 58124 26732 58130 26744
rect 58253 26741 58265 26744
rect 58299 26741 58311 26775
rect 58253 26735 58311 26741
rect 1104 26682 68816 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 68816 26682
rect 1104 26608 68816 26630
rect 33778 26568 33784 26580
rect 33739 26540 33784 26568
rect 33778 26528 33784 26540
rect 33836 26528 33842 26580
rect 34790 26568 34796 26580
rect 34751 26540 34796 26568
rect 34790 26528 34796 26540
rect 34848 26528 34854 26580
rect 55766 26432 55772 26444
rect 55727 26404 55772 26432
rect 55766 26392 55772 26404
rect 55824 26392 55830 26444
rect 58066 26432 58072 26444
rect 58027 26404 58072 26432
rect 58066 26392 58072 26404
rect 58124 26392 58130 26444
rect 26145 26367 26203 26373
rect 26145 26333 26157 26367
rect 26191 26364 26203 26367
rect 26878 26364 26884 26376
rect 26191 26336 26884 26364
rect 26191 26333 26203 26336
rect 26145 26327 26203 26333
rect 26878 26324 26884 26336
rect 26936 26324 26942 26376
rect 34885 26367 34943 26373
rect 34885 26333 34897 26367
rect 34931 26364 34943 26367
rect 35342 26364 35348 26376
rect 34931 26336 35348 26364
rect 34931 26333 34943 26336
rect 34885 26327 34943 26333
rect 35342 26324 35348 26336
rect 35400 26324 35406 26376
rect 59909 26367 59967 26373
rect 59909 26333 59921 26367
rect 59955 26364 59967 26367
rect 66162 26364 66168 26376
rect 59955 26336 66168 26364
rect 59955 26333 59967 26336
rect 59909 26327 59967 26333
rect 66162 26324 66168 26336
rect 66220 26324 66226 26376
rect 55950 26296 55956 26308
rect 55911 26268 55956 26296
rect 55950 26256 55956 26268
rect 56008 26256 56014 26308
rect 57606 26296 57612 26308
rect 57567 26268 57612 26296
rect 57606 26256 57612 26268
rect 57664 26256 57670 26308
rect 58250 26296 58256 26308
rect 58211 26268 58256 26296
rect 58250 26256 58256 26268
rect 58308 26256 58314 26308
rect 1104 26138 68816 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 68816 26138
rect 1104 26064 68816 26086
rect 55950 25984 55956 26036
rect 56008 26024 56014 26036
rect 56413 26027 56471 26033
rect 56413 26024 56425 26027
rect 56008 25996 56425 26024
rect 56008 25984 56014 25996
rect 56413 25993 56425 25996
rect 56459 25993 56471 26027
rect 58250 26024 58256 26036
rect 58211 25996 58256 26024
rect 56413 25987 56471 25993
rect 58250 25984 58256 25996
rect 58308 25984 58314 26036
rect 27154 25888 27160 25900
rect 27115 25860 27160 25888
rect 27154 25848 27160 25860
rect 27212 25848 27218 25900
rect 56502 25888 56508 25900
rect 56463 25860 56508 25888
rect 56502 25848 56508 25860
rect 56560 25848 56566 25900
rect 58158 25888 58164 25900
rect 58119 25860 58164 25888
rect 58158 25848 58164 25860
rect 58216 25848 58222 25900
rect 27065 25687 27123 25693
rect 27065 25653 27077 25687
rect 27111 25684 27123 25687
rect 27522 25684 27528 25696
rect 27111 25656 27528 25684
rect 27111 25653 27123 25656
rect 27065 25647 27123 25653
rect 27522 25644 27528 25656
rect 27580 25644 27586 25696
rect 1104 25594 68816 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 68816 25594
rect 1104 25520 68816 25542
rect 26878 25372 26884 25424
rect 26936 25412 26942 25424
rect 26936 25384 27752 25412
rect 26936 25372 26942 25384
rect 27522 25344 27528 25356
rect 27483 25316 27528 25344
rect 27522 25304 27528 25316
rect 27580 25304 27586 25356
rect 27724 25353 27752 25384
rect 27709 25347 27767 25353
rect 27709 25313 27721 25347
rect 27755 25313 27767 25347
rect 27709 25307 27767 25313
rect 32122 25304 32128 25356
rect 32180 25344 32186 25356
rect 32677 25347 32735 25353
rect 32677 25344 32689 25347
rect 32180 25316 32689 25344
rect 32180 25304 32186 25316
rect 32677 25313 32689 25316
rect 32723 25313 32735 25347
rect 32677 25307 32735 25313
rect 12342 25276 12348 25288
rect 12303 25248 12348 25276
rect 12342 25236 12348 25248
rect 12400 25236 12406 25288
rect 28166 25276 28172 25288
rect 28127 25248 28172 25276
rect 28166 25236 28172 25248
rect 28224 25236 28230 25288
rect 32217 25279 32275 25285
rect 32217 25245 32229 25279
rect 32263 25276 32275 25279
rect 35710 25276 35716 25288
rect 32263 25248 35716 25276
rect 32263 25245 32275 25248
rect 32217 25239 32275 25245
rect 35710 25236 35716 25248
rect 35768 25236 35774 25288
rect 3142 25168 3148 25220
rect 3200 25208 3206 25220
rect 25869 25211 25927 25217
rect 25869 25208 25881 25211
rect 3200 25180 25881 25208
rect 3200 25168 3206 25180
rect 25869 25177 25881 25180
rect 25915 25177 25927 25211
rect 25869 25171 25927 25177
rect 32125 25143 32183 25149
rect 32125 25109 32137 25143
rect 32171 25140 32183 25143
rect 32306 25140 32312 25152
rect 32171 25112 32312 25140
rect 32171 25109 32183 25112
rect 32125 25103 32183 25109
rect 32306 25100 32312 25112
rect 32364 25100 32370 25152
rect 1104 25050 68816 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 68816 25050
rect 1104 24976 68816 24998
rect 27154 24896 27160 24948
rect 27212 24936 27218 24948
rect 33686 24936 33692 24948
rect 27212 24908 33692 24936
rect 27212 24896 27218 24908
rect 33686 24896 33692 24908
rect 33744 24896 33750 24948
rect 32306 24868 32312 24880
rect 32267 24840 32312 24868
rect 32306 24828 32312 24840
rect 32364 24828 32370 24880
rect 12342 24800 12348 24812
rect 12303 24772 12348 24800
rect 12342 24760 12348 24772
rect 12400 24760 12406 24812
rect 23661 24803 23719 24809
rect 23661 24769 23673 24803
rect 23707 24800 23719 24803
rect 27982 24800 27988 24812
rect 23707 24772 27988 24800
rect 23707 24769 23719 24772
rect 23661 24763 23719 24769
rect 27982 24760 27988 24772
rect 28040 24760 28046 24812
rect 28166 24800 28172 24812
rect 28127 24772 28172 24800
rect 28166 24760 28172 24772
rect 28224 24760 28230 24812
rect 32122 24800 32128 24812
rect 32083 24772 32128 24800
rect 32122 24760 32128 24772
rect 32180 24760 32186 24812
rect 12529 24735 12587 24741
rect 12529 24701 12541 24735
rect 12575 24732 12587 24735
rect 12986 24732 12992 24744
rect 12575 24704 12992 24732
rect 12575 24701 12587 24704
rect 12529 24695 12587 24701
rect 12986 24692 12992 24704
rect 13044 24692 13050 24744
rect 13081 24735 13139 24741
rect 13081 24701 13093 24735
rect 13127 24701 13139 24735
rect 13081 24695 13139 24701
rect 28353 24735 28411 24741
rect 28353 24701 28365 24735
rect 28399 24732 28411 24735
rect 28534 24732 28540 24744
rect 28399 24704 28540 24732
rect 28399 24701 28411 24704
rect 28353 24695 28411 24701
rect 3418 24624 3424 24676
rect 3476 24664 3482 24676
rect 13096 24664 13124 24695
rect 28534 24692 28540 24704
rect 28592 24692 28598 24744
rect 28629 24735 28687 24741
rect 28629 24701 28641 24735
rect 28675 24701 28687 24735
rect 28629 24695 28687 24701
rect 32585 24735 32643 24741
rect 32585 24701 32597 24735
rect 32631 24701 32643 24735
rect 32585 24695 32643 24701
rect 28644 24664 28672 24695
rect 3476 24636 13124 24664
rect 16546 24636 28672 24664
rect 3476 24624 3482 24636
rect 3602 24556 3608 24608
rect 3660 24596 3666 24608
rect 16546 24596 16574 24636
rect 31754 24624 31760 24676
rect 31812 24664 31818 24676
rect 32600 24664 32628 24695
rect 31812 24636 32628 24664
rect 31812 24624 31818 24636
rect 23014 24596 23020 24608
rect 3660 24568 16574 24596
rect 22975 24568 23020 24596
rect 3660 24556 3666 24568
rect 23014 24556 23020 24568
rect 23072 24556 23078 24608
rect 23198 24556 23204 24608
rect 23256 24596 23262 24608
rect 23569 24599 23627 24605
rect 23569 24596 23581 24599
rect 23256 24568 23581 24596
rect 23256 24556 23262 24568
rect 23569 24565 23581 24568
rect 23615 24565 23627 24599
rect 23569 24559 23627 24565
rect 27982 24556 27988 24608
rect 28040 24596 28046 24608
rect 35434 24596 35440 24608
rect 28040 24568 35440 24596
rect 28040 24556 28046 24568
rect 35434 24556 35440 24568
rect 35492 24556 35498 24608
rect 1104 24506 68816 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 68816 24506
rect 1104 24432 68816 24454
rect 12986 24392 12992 24404
rect 12947 24364 12992 24392
rect 12986 24352 12992 24364
rect 13044 24352 13050 24404
rect 28534 24392 28540 24404
rect 28495 24364 28540 24392
rect 28534 24352 28540 24364
rect 28592 24352 28598 24404
rect 13081 24191 13139 24197
rect 13081 24157 13093 24191
rect 13127 24188 13139 24191
rect 14274 24188 14280 24200
rect 13127 24160 14280 24188
rect 13127 24157 13139 24160
rect 13081 24151 13139 24157
rect 14274 24148 14280 24160
rect 14332 24188 14338 24200
rect 14458 24188 14464 24200
rect 14332 24160 14464 24188
rect 14332 24148 14338 24160
rect 14458 24148 14464 24160
rect 14516 24148 14522 24200
rect 28629 24191 28687 24197
rect 28629 24157 28641 24191
rect 28675 24188 28687 24191
rect 34790 24188 34796 24200
rect 28675 24160 34796 24188
rect 28675 24157 28687 24160
rect 28629 24151 28687 24157
rect 34790 24148 34796 24160
rect 34848 24148 34854 24200
rect 1104 23962 68816 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 68816 23962
rect 1104 23888 68816 23910
rect 23198 23780 23204 23792
rect 23159 23752 23204 23780
rect 23198 23740 23204 23752
rect 23256 23740 23262 23792
rect 23014 23712 23020 23724
rect 22975 23684 23020 23712
rect 23014 23672 23020 23684
rect 23072 23672 23078 23724
rect 24670 23644 24676 23656
rect 24631 23616 24676 23644
rect 24670 23604 24676 23616
rect 24728 23604 24734 23656
rect 1104 23418 68816 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 68816 23418
rect 1104 23344 68816 23366
rect 1104 22874 68816 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 68816 22874
rect 1104 22800 68816 22822
rect 51721 22695 51779 22701
rect 51721 22661 51733 22695
rect 51767 22692 51779 22695
rect 52917 22695 52975 22701
rect 52917 22692 52929 22695
rect 51767 22664 52929 22692
rect 51767 22661 51779 22664
rect 51721 22655 51779 22661
rect 52917 22661 52929 22664
rect 52963 22661 52975 22695
rect 52917 22655 52975 22661
rect 35342 22584 35348 22636
rect 35400 22624 35406 22636
rect 51629 22627 51687 22633
rect 51629 22624 51641 22627
rect 35400 22596 51641 22624
rect 35400 22584 35406 22596
rect 51629 22593 51641 22596
rect 51675 22593 51687 22627
rect 51629 22587 51687 22593
rect 52178 22516 52184 22568
rect 52236 22556 52242 22568
rect 52733 22559 52791 22565
rect 52733 22556 52745 22559
rect 52236 22528 52745 22556
rect 52236 22516 52242 22528
rect 52733 22525 52745 22528
rect 52779 22525 52791 22559
rect 54570 22556 54576 22568
rect 54531 22528 54576 22556
rect 52733 22519 52791 22525
rect 54570 22516 54576 22528
rect 54628 22516 54634 22568
rect 6549 22423 6607 22429
rect 6549 22389 6561 22423
rect 6595 22420 6607 22423
rect 7558 22420 7564 22432
rect 6595 22392 7564 22420
rect 6595 22389 6607 22392
rect 6549 22383 6607 22389
rect 7558 22380 7564 22392
rect 7616 22380 7622 22432
rect 9306 22420 9312 22432
rect 9267 22392 9312 22420
rect 9306 22380 9312 22392
rect 9364 22380 9370 22432
rect 11698 22380 11704 22432
rect 11756 22420 11762 22432
rect 11793 22423 11851 22429
rect 11793 22420 11805 22423
rect 11756 22392 11805 22420
rect 11756 22380 11762 22392
rect 11793 22389 11805 22392
rect 11839 22389 11851 22423
rect 11793 22383 11851 22389
rect 56318 22380 56324 22432
rect 56376 22420 56382 22432
rect 56413 22423 56471 22429
rect 56413 22420 56425 22423
rect 56376 22392 56425 22420
rect 56376 22380 56382 22392
rect 56413 22389 56425 22392
rect 56459 22389 56471 22423
rect 56413 22383 56471 22389
rect 61746 22380 61752 22432
rect 61804 22420 61810 22432
rect 61841 22423 61899 22429
rect 61841 22420 61853 22423
rect 61804 22392 61853 22420
rect 61804 22380 61810 22392
rect 61841 22389 61853 22392
rect 61887 22389 61899 22423
rect 61841 22383 61899 22389
rect 1104 22330 68816 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 68816 22330
rect 1104 22256 68816 22278
rect 52178 22216 52184 22228
rect 52139 22188 52184 22216
rect 52178 22176 52184 22188
rect 52236 22176 52242 22228
rect 7392 22120 7696 22148
rect 3510 22040 3516 22092
rect 3568 22080 3574 22092
rect 7392 22080 7420 22120
rect 7558 22080 7564 22092
rect 3568 22052 7420 22080
rect 7519 22052 7564 22080
rect 3568 22040 3574 22052
rect 7558 22040 7564 22052
rect 7616 22040 7622 22092
rect 4614 21904 4620 21956
rect 4672 21944 4678 21956
rect 5721 21947 5779 21953
rect 5721 21944 5733 21947
rect 4672 21916 5733 21944
rect 4672 21904 4678 21916
rect 5721 21913 5733 21916
rect 5767 21913 5779 21947
rect 5721 21907 5779 21913
rect 6454 21904 6460 21956
rect 6512 21944 6518 21956
rect 7377 21947 7435 21953
rect 7377 21944 7389 21947
rect 6512 21916 7389 21944
rect 6512 21904 6518 21916
rect 7377 21913 7389 21916
rect 7423 21913 7435 21947
rect 7668 21944 7696 22120
rect 26436 22120 26740 22148
rect 9306 22080 9312 22092
rect 9267 22052 9312 22080
rect 9306 22040 9312 22052
rect 9364 22040 9370 22092
rect 9490 22080 9496 22092
rect 9451 22052 9496 22080
rect 9490 22040 9496 22052
rect 9548 22040 9554 22092
rect 9766 22080 9772 22092
rect 9727 22052 9772 22080
rect 9766 22040 9772 22052
rect 9824 22040 9830 22092
rect 11698 22080 11704 22092
rect 11659 22052 11704 22080
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 13081 22083 13139 22089
rect 13081 22049 13093 22083
rect 13127 22049 13139 22083
rect 26436 22080 26464 22120
rect 26602 22080 26608 22092
rect 13081 22043 13139 22049
rect 25516 22052 26464 22080
rect 26563 22052 26608 22080
rect 11885 21947 11943 21953
rect 7668 21916 9996 21944
rect 7377 21907 7435 21913
rect 4062 21836 4068 21888
rect 4120 21876 4126 21888
rect 9766 21876 9772 21888
rect 4120 21848 9772 21876
rect 4120 21836 4126 21848
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 9968 21876 9996 21916
rect 11885 21913 11897 21947
rect 11931 21944 11943 21947
rect 12066 21944 12072 21956
rect 11931 21916 12072 21944
rect 11931 21913 11943 21916
rect 11885 21907 11943 21913
rect 12066 21904 12072 21916
rect 12124 21904 12130 21956
rect 13096 21876 13124 22043
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 25516 22021 25544 22052
rect 26602 22040 26608 22052
rect 26660 22040 26666 22092
rect 26712 22080 26740 22120
rect 35526 22080 35532 22092
rect 26712 22052 35532 22080
rect 35526 22040 35532 22052
rect 35584 22040 35590 22092
rect 56318 22080 56324 22092
rect 56279 22052 56324 22080
rect 56318 22040 56324 22052
rect 56376 22040 56382 22092
rect 57882 22080 57888 22092
rect 57843 22052 57888 22080
rect 57882 22040 57888 22052
rect 57940 22040 57946 22092
rect 61746 22080 61752 22092
rect 61707 22052 61752 22080
rect 61746 22040 61752 22052
rect 61804 22040 61810 22092
rect 25501 22015 25559 22021
rect 25501 22012 25513 22015
rect 24820 21984 25513 22012
rect 24820 21972 24826 21984
rect 25501 21981 25513 21984
rect 25547 21981 25559 22015
rect 26142 22012 26148 22024
rect 26103 21984 26148 22012
rect 25501 21975 25559 21981
rect 26142 21972 26148 21984
rect 26200 21972 26206 22024
rect 25593 21947 25651 21953
rect 25593 21913 25605 21947
rect 25639 21944 25651 21947
rect 26329 21947 26387 21953
rect 26329 21944 26341 21947
rect 25639 21916 26341 21944
rect 25639 21913 25651 21916
rect 25593 21907 25651 21913
rect 26329 21913 26341 21916
rect 26375 21913 26387 21947
rect 26329 21907 26387 21913
rect 56318 21904 56324 21956
rect 56376 21944 56382 21956
rect 56505 21947 56563 21953
rect 56505 21944 56517 21947
rect 56376 21916 56517 21944
rect 56376 21904 56382 21916
rect 56505 21913 56517 21916
rect 56551 21913 56563 21947
rect 56505 21907 56563 21913
rect 61746 21904 61752 21956
rect 61804 21944 61810 21956
rect 61933 21947 61991 21953
rect 61933 21944 61945 21947
rect 61804 21916 61945 21944
rect 61804 21904 61810 21916
rect 61933 21913 61945 21916
rect 61979 21913 61991 21947
rect 61933 21907 61991 21913
rect 63589 21947 63647 21953
rect 63589 21913 63601 21947
rect 63635 21944 63647 21947
rect 66162 21944 66168 21956
rect 63635 21916 66168 21944
rect 63635 21913 63647 21916
rect 63589 21907 63647 21913
rect 66162 21904 66168 21916
rect 66220 21904 66226 21956
rect 9968 21848 13124 21876
rect 1104 21786 68816 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 68816 21786
rect 1104 21712 68816 21734
rect 6454 21672 6460 21684
rect 6415 21644 6460 21672
rect 6454 21632 6460 21644
rect 6512 21632 6518 21684
rect 9490 21632 9496 21684
rect 9548 21672 9554 21684
rect 9677 21675 9735 21681
rect 9677 21672 9689 21675
rect 9548 21644 9689 21672
rect 9548 21632 9554 21644
rect 9677 21641 9689 21644
rect 9723 21641 9735 21675
rect 12066 21672 12072 21684
rect 12027 21644 12072 21672
rect 9677 21635 9735 21641
rect 12066 21632 12072 21644
rect 12124 21632 12130 21684
rect 26602 21672 26608 21684
rect 16546 21644 26608 21672
rect 9784 21576 12296 21604
rect 6546 21536 6552 21548
rect 6507 21508 6552 21536
rect 6546 21496 6552 21508
rect 6604 21496 6610 21548
rect 9674 21496 9680 21548
rect 9732 21536 9738 21548
rect 9784 21545 9812 21576
rect 9769 21539 9827 21545
rect 9769 21536 9781 21539
rect 9732 21508 9781 21536
rect 9732 21496 9738 21508
rect 9769 21505 9781 21508
rect 9815 21505 9827 21539
rect 9769 21499 9827 21505
rect 11790 21496 11796 21548
rect 11848 21536 11854 21548
rect 12161 21539 12219 21545
rect 12161 21536 12173 21539
rect 11848 21508 12173 21536
rect 11848 21496 11854 21508
rect 12161 21505 12173 21508
rect 12207 21505 12219 21539
rect 12268 21536 12296 21576
rect 12342 21564 12348 21616
rect 12400 21604 12406 21616
rect 16546 21604 16574 21644
rect 26602 21632 26608 21644
rect 26660 21632 26666 21684
rect 56318 21672 56324 21684
rect 56279 21644 56324 21672
rect 56318 21632 56324 21644
rect 56376 21632 56382 21684
rect 61746 21672 61752 21684
rect 61707 21644 61752 21672
rect 61746 21632 61752 21644
rect 61804 21632 61810 21684
rect 12400 21576 16574 21604
rect 12400 21564 12406 21576
rect 36446 21536 36452 21548
rect 12268 21508 36452 21536
rect 12161 21499 12219 21505
rect 12176 21332 12204 21499
rect 36446 21496 36452 21508
rect 36504 21496 36510 21548
rect 56229 21539 56287 21545
rect 56229 21505 56241 21539
rect 56275 21536 56287 21539
rect 56502 21536 56508 21548
rect 56275 21508 56508 21536
rect 56275 21505 56287 21508
rect 56229 21499 56287 21505
rect 56502 21496 56508 21508
rect 56560 21496 56566 21548
rect 61654 21536 61660 21548
rect 61615 21508 61660 21536
rect 61654 21496 61660 21508
rect 61712 21496 61718 21548
rect 17862 21468 17868 21480
rect 16546 21440 17868 21468
rect 16546 21332 16574 21440
rect 17862 21428 17868 21440
rect 17920 21428 17926 21480
rect 26142 21428 26148 21480
rect 26200 21468 26206 21480
rect 26237 21471 26295 21477
rect 26237 21468 26249 21471
rect 26200 21440 26249 21468
rect 26200 21428 26206 21440
rect 26237 21437 26249 21440
rect 26283 21437 26295 21471
rect 26237 21431 26295 21437
rect 12176 21304 16574 21332
rect 1104 21242 68816 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 68816 21242
rect 1104 21168 68816 21190
rect 3970 21088 3976 21140
rect 4028 21128 4034 21140
rect 12342 21128 12348 21140
rect 4028 21100 12348 21128
rect 4028 21088 4034 21100
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 17862 20952 17868 21004
rect 17920 20992 17926 21004
rect 27341 20995 27399 21001
rect 27341 20992 27353 20995
rect 17920 20964 27353 20992
rect 17920 20952 17926 20964
rect 27341 20961 27353 20964
rect 27387 20961 27399 20995
rect 27341 20955 27399 20961
rect 8662 20884 8668 20936
rect 8720 20924 8726 20936
rect 8941 20927 8999 20933
rect 8941 20924 8953 20927
rect 8720 20896 8953 20924
rect 8720 20884 8726 20896
rect 8941 20893 8953 20896
rect 8987 20893 8999 20927
rect 27154 20924 27160 20936
rect 27115 20896 27160 20924
rect 8941 20887 8999 20893
rect 27154 20884 27160 20896
rect 27212 20884 27218 20936
rect 62666 20924 62672 20936
rect 62627 20896 62672 20924
rect 62666 20884 62672 20896
rect 62724 20884 62730 20936
rect 1104 20698 68816 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 68816 20698
rect 1104 20624 68816 20646
rect 8662 20448 8668 20460
rect 8623 20420 8668 20448
rect 8662 20408 8668 20420
rect 8720 20408 8726 20460
rect 61654 20408 61660 20460
rect 61712 20448 61718 20460
rect 62022 20448 62028 20460
rect 61712 20420 62028 20448
rect 61712 20408 61718 20420
rect 62022 20408 62028 20420
rect 62080 20448 62086 20460
rect 62209 20451 62267 20457
rect 62209 20448 62221 20451
rect 62080 20420 62221 20448
rect 62080 20408 62086 20420
rect 62209 20417 62221 20420
rect 62255 20417 62267 20451
rect 62209 20411 62267 20417
rect 62666 20408 62672 20460
rect 62724 20448 62730 20460
rect 63037 20451 63095 20457
rect 63037 20448 63049 20451
rect 62724 20420 63049 20448
rect 62724 20408 62730 20420
rect 63037 20417 63049 20420
rect 63083 20417 63095 20451
rect 63037 20411 63095 20417
rect 64874 20408 64880 20460
rect 64932 20448 64938 20460
rect 64932 20420 64977 20448
rect 64932 20408 64938 20420
rect 8849 20383 8907 20389
rect 8849 20349 8861 20383
rect 8895 20380 8907 20383
rect 9030 20380 9036 20392
rect 8895 20352 9036 20380
rect 8895 20349 8907 20352
rect 8849 20343 8907 20349
rect 9030 20340 9036 20352
rect 9088 20340 9094 20392
rect 9125 20383 9183 20389
rect 9125 20349 9137 20383
rect 9171 20349 9183 20383
rect 9125 20343 9183 20349
rect 62301 20383 62359 20389
rect 62301 20349 62313 20383
rect 62347 20380 62359 20383
rect 63221 20383 63279 20389
rect 63221 20380 63233 20383
rect 62347 20352 63233 20380
rect 62347 20349 62359 20352
rect 62301 20343 62359 20349
rect 63221 20349 63233 20352
rect 63267 20349 63279 20383
rect 63221 20343 63279 20349
rect 4062 20272 4068 20324
rect 4120 20312 4126 20324
rect 9140 20312 9168 20343
rect 4120 20284 9168 20312
rect 4120 20272 4126 20284
rect 1104 20154 68816 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 68816 20154
rect 1104 20080 68816 20102
rect 9030 20040 9036 20052
rect 8991 20012 9036 20040
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 8386 19796 8392 19848
rect 8444 19836 8450 19848
rect 9122 19836 9128 19848
rect 8444 19808 9128 19836
rect 8444 19796 8450 19808
rect 9122 19796 9128 19808
rect 9180 19796 9186 19848
rect 1104 19610 68816 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 68816 19610
rect 1104 19536 68816 19558
rect 27890 19360 27896 19372
rect 27851 19332 27896 19360
rect 27890 19320 27896 19332
rect 27948 19320 27954 19372
rect 34698 19320 34704 19372
rect 34756 19360 34762 19372
rect 35161 19363 35219 19369
rect 35161 19360 35173 19363
rect 34756 19332 35173 19360
rect 34756 19320 34762 19332
rect 35161 19329 35173 19332
rect 35207 19329 35219 19363
rect 35161 19323 35219 19329
rect 53374 19252 53380 19304
rect 53432 19292 53438 19304
rect 66162 19292 66168 19304
rect 53432 19264 66168 19292
rect 53432 19252 53438 19264
rect 66162 19252 66168 19264
rect 66220 19252 66226 19304
rect 35253 19227 35311 19233
rect 35253 19193 35265 19227
rect 35299 19224 35311 19227
rect 35710 19224 35716 19236
rect 35299 19196 35716 19224
rect 35299 19193 35311 19196
rect 35253 19187 35311 19193
rect 35710 19184 35716 19196
rect 35768 19184 35774 19236
rect 27982 19156 27988 19168
rect 27943 19128 27988 19156
rect 27982 19116 27988 19128
rect 28040 19116 28046 19168
rect 28721 19159 28779 19165
rect 28721 19125 28733 19159
rect 28767 19156 28779 19159
rect 28994 19156 29000 19168
rect 28767 19128 29000 19156
rect 28767 19125 28779 19128
rect 28721 19119 28779 19125
rect 28994 19116 29000 19128
rect 29052 19116 29058 19168
rect 35526 19116 35532 19168
rect 35584 19156 35590 19168
rect 35805 19159 35863 19165
rect 35805 19156 35817 19159
rect 35584 19128 35817 19156
rect 35584 19116 35590 19128
rect 35805 19125 35817 19128
rect 35851 19125 35863 19159
rect 35805 19119 35863 19125
rect 1104 19066 68816 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 68816 19066
rect 1104 18992 68816 19014
rect 27982 18776 27988 18828
rect 28040 18816 28046 18828
rect 28813 18819 28871 18825
rect 28813 18816 28825 18819
rect 28040 18788 28825 18816
rect 28040 18776 28046 18788
rect 28813 18785 28825 18788
rect 28859 18785 28871 18819
rect 28994 18816 29000 18828
rect 28955 18788 29000 18816
rect 28813 18779 28871 18785
rect 28994 18776 29000 18788
rect 29052 18776 29058 18828
rect 35526 18816 35532 18828
rect 35487 18788 35532 18816
rect 35526 18776 35532 18788
rect 35584 18776 35590 18828
rect 35710 18816 35716 18828
rect 35671 18788 35716 18816
rect 35710 18776 35716 18788
rect 35768 18776 35774 18828
rect 37182 18816 37188 18828
rect 37143 18788 37188 18816
rect 37182 18776 37188 18788
rect 37240 18776 37246 18828
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18748 23903 18751
rect 24118 18748 24124 18760
rect 23891 18720 24124 18748
rect 23891 18717 23903 18720
rect 23845 18711 23903 18717
rect 24118 18708 24124 18720
rect 24176 18708 24182 18760
rect 24762 18748 24768 18760
rect 24723 18720 24768 18748
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 4706 18640 4712 18692
rect 4764 18680 4770 18692
rect 27157 18683 27215 18689
rect 27157 18680 27169 18683
rect 4764 18652 27169 18680
rect 4764 18640 4770 18652
rect 27157 18649 27169 18652
rect 27203 18649 27215 18683
rect 27157 18643 27215 18649
rect 24302 18572 24308 18624
rect 24360 18612 24366 18624
rect 24673 18615 24731 18621
rect 24673 18612 24685 18615
rect 24360 18584 24685 18612
rect 24360 18572 24366 18584
rect 24673 18581 24685 18584
rect 24719 18581 24731 18615
rect 24673 18575 24731 18581
rect 1104 18522 68816 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 68816 18522
rect 1104 18448 68816 18470
rect 24302 18340 24308 18352
rect 24263 18312 24308 18340
rect 24302 18300 24308 18312
rect 24360 18300 24366 18352
rect 24118 18272 24124 18284
rect 24079 18244 24124 18272
rect 24118 18232 24124 18244
rect 24176 18232 24182 18284
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 24136 18176 24593 18204
rect 24136 18148 24164 18176
rect 24581 18173 24593 18176
rect 24627 18173 24639 18207
rect 24581 18167 24639 18173
rect 24118 18096 24124 18148
rect 24176 18096 24182 18148
rect 1104 17978 68816 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 68816 17978
rect 1104 17904 68816 17926
rect 52914 17824 52920 17876
rect 52972 17864 52978 17876
rect 66162 17864 66168 17876
rect 52972 17836 66168 17864
rect 52972 17824 52978 17836
rect 66162 17824 66168 17836
rect 66220 17824 66226 17876
rect 38470 17728 38476 17740
rect 38431 17700 38476 17728
rect 38470 17688 38476 17700
rect 38528 17688 38534 17740
rect 13722 17620 13728 17672
rect 13780 17660 13786 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13780 17632 14105 17660
rect 13780 17620 13786 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 33686 17620 33692 17672
rect 33744 17660 33750 17672
rect 36173 17663 36231 17669
rect 36173 17660 36185 17663
rect 33744 17632 36185 17660
rect 33744 17620 33750 17632
rect 36173 17629 36185 17632
rect 36219 17629 36231 17663
rect 36814 17660 36820 17672
rect 36775 17632 36820 17660
rect 36173 17623 36231 17629
rect 36814 17620 36820 17632
rect 36872 17620 36878 17672
rect 58158 17620 58164 17672
rect 58216 17660 58222 17672
rect 58805 17663 58863 17669
rect 58805 17660 58817 17663
rect 58216 17632 58817 17660
rect 58216 17620 58222 17632
rect 58805 17629 58817 17632
rect 58851 17629 58863 17663
rect 58805 17623 58863 17629
rect 59170 17620 59176 17672
rect 59228 17660 59234 17672
rect 59449 17663 59507 17669
rect 59449 17660 59461 17663
rect 59228 17632 59461 17660
rect 59228 17620 59234 17632
rect 59449 17629 59461 17632
rect 59495 17629 59507 17663
rect 59449 17623 59507 17629
rect 36265 17595 36323 17601
rect 36265 17561 36277 17595
rect 36311 17592 36323 17595
rect 37001 17595 37059 17601
rect 37001 17592 37013 17595
rect 36311 17564 37013 17592
rect 36311 17561 36323 17564
rect 36265 17555 36323 17561
rect 37001 17561 37013 17564
rect 37047 17561 37059 17595
rect 37001 17555 37059 17561
rect 58897 17527 58955 17533
rect 58897 17493 58909 17527
rect 58943 17524 58955 17527
rect 59354 17524 59360 17536
rect 58943 17496 59360 17524
rect 58943 17493 58955 17496
rect 58897 17487 58955 17493
rect 59354 17484 59360 17496
rect 59412 17484 59418 17536
rect 1104 17434 68816 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 68816 17434
rect 1104 17360 68816 17382
rect 59354 17252 59360 17264
rect 59315 17224 59360 17252
rect 59354 17212 59360 17224
rect 59412 17212 59418 17264
rect 13722 17184 13728 17196
rect 13683 17156 13728 17184
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 36814 17144 36820 17196
rect 36872 17184 36878 17196
rect 37277 17187 37335 17193
rect 37277 17184 37289 17187
rect 36872 17156 37289 17184
rect 36872 17144 36878 17156
rect 37277 17153 37289 17156
rect 37323 17153 37335 17187
rect 59170 17184 59176 17196
rect 59131 17156 59176 17184
rect 37277 17147 37335 17153
rect 59170 17144 59176 17156
rect 59228 17144 59234 17196
rect 13906 17116 13912 17128
rect 13867 17088 13912 17116
rect 13906 17076 13912 17088
rect 13964 17076 13970 17128
rect 14458 17116 14464 17128
rect 14419 17088 14464 17116
rect 14458 17076 14464 17088
rect 14516 17076 14522 17128
rect 61013 17119 61071 17125
rect 61013 17085 61025 17119
rect 61059 17116 61071 17119
rect 65518 17116 65524 17128
rect 61059 17088 65524 17116
rect 61059 17085 61071 17088
rect 61013 17079 61071 17085
rect 65518 17076 65524 17088
rect 65576 17076 65582 17128
rect 1104 16890 68816 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 68816 16890
rect 1104 16816 68816 16838
rect 13906 16736 13912 16788
rect 13964 16776 13970 16788
rect 14185 16779 14243 16785
rect 14185 16776 14197 16779
rect 13964 16748 14197 16776
rect 13964 16736 13970 16748
rect 14185 16745 14197 16748
rect 14231 16745 14243 16779
rect 14185 16739 14243 16745
rect 14274 16582 14280 16594
rect 14235 16554 14280 16582
rect 14274 16542 14280 16554
rect 14332 16542 14338 16594
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 4614 16436 4620 16448
rect 4120 16408 4620 16436
rect 4120 16396 4126 16408
rect 4614 16396 4620 16408
rect 4672 16396 4678 16448
rect 1104 16346 68816 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 68816 16346
rect 1104 16272 68816 16294
rect 1104 15802 68816 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 68816 15802
rect 1104 15728 68816 15750
rect 23106 15444 23112 15496
rect 23164 15484 23170 15496
rect 23201 15487 23259 15493
rect 23201 15484 23213 15487
rect 23164 15456 23213 15484
rect 23164 15444 23170 15456
rect 23201 15453 23213 15456
rect 23247 15453 23259 15487
rect 23201 15447 23259 15453
rect 23845 15487 23903 15493
rect 23845 15453 23857 15487
rect 23891 15484 23903 15487
rect 27890 15484 27896 15496
rect 23891 15456 27896 15484
rect 23891 15453 23903 15456
rect 23845 15447 23903 15453
rect 27890 15444 27896 15456
rect 27948 15444 27954 15496
rect 62022 15484 62028 15496
rect 61983 15456 62028 15484
rect 62022 15444 62028 15456
rect 62080 15444 62086 15496
rect 62850 15484 62856 15496
rect 62811 15456 62856 15484
rect 62850 15444 62856 15456
rect 62908 15444 62914 15496
rect 23750 15348 23756 15360
rect 23711 15320 23756 15348
rect 23750 15308 23756 15320
rect 23808 15308 23814 15360
rect 62117 15351 62175 15357
rect 62117 15317 62129 15351
rect 62163 15348 62175 15351
rect 63218 15348 63224 15360
rect 62163 15320 63224 15348
rect 62163 15317 62175 15320
rect 62117 15311 62175 15317
rect 63218 15308 63224 15320
rect 63276 15308 63282 15360
rect 1104 15258 68816 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 68816 15258
rect 1104 15184 68816 15206
rect 23293 15079 23351 15085
rect 23293 15045 23305 15079
rect 23339 15076 23351 15079
rect 23750 15076 23756 15088
rect 23339 15048 23756 15076
rect 23339 15045 23351 15048
rect 23293 15039 23351 15045
rect 23750 15036 23756 15048
rect 23808 15036 23814 15088
rect 63218 15076 63224 15088
rect 63179 15048 63224 15076
rect 63218 15036 63224 15048
rect 63276 15036 63282 15088
rect 23106 15008 23112 15020
rect 23067 14980 23112 15008
rect 23106 14968 23112 14980
rect 23164 14968 23170 15020
rect 62850 14968 62856 15020
rect 62908 15008 62914 15020
rect 63037 15011 63095 15017
rect 63037 15008 63049 15011
rect 62908 14980 63049 15008
rect 62908 14968 62914 14980
rect 63037 14977 63049 14980
rect 63083 14977 63095 15011
rect 63037 14971 63095 14977
rect 23569 14943 23627 14949
rect 23569 14940 23581 14943
rect 2746 14912 23581 14940
rect 842 14832 848 14884
rect 900 14872 906 14884
rect 2746 14872 2774 14912
rect 23569 14909 23581 14912
rect 23615 14909 23627 14943
rect 64782 14940 64788 14952
rect 64743 14912 64788 14940
rect 23569 14903 23627 14909
rect 64782 14900 64788 14912
rect 64840 14900 64846 14952
rect 900 14844 2774 14872
rect 900 14832 906 14844
rect 1104 14714 68816 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 68816 14714
rect 1104 14640 68816 14662
rect 38838 14464 38844 14476
rect 35866 14436 38844 14464
rect 14274 14356 14280 14408
rect 14332 14396 14338 14408
rect 15013 14399 15071 14405
rect 15013 14396 15025 14399
rect 14332 14368 15025 14396
rect 14332 14356 14338 14368
rect 15013 14365 15025 14368
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 35713 14399 35771 14405
rect 35713 14365 35725 14399
rect 35759 14396 35771 14399
rect 35866 14396 35894 14436
rect 38838 14424 38844 14436
rect 38896 14424 38902 14476
rect 36354 14396 36360 14408
rect 35759 14368 35894 14396
rect 36315 14368 36360 14396
rect 35759 14365 35771 14368
rect 35713 14359 35771 14365
rect 36354 14356 36360 14368
rect 36412 14356 36418 14408
rect 15102 14260 15108 14272
rect 15063 14232 15108 14260
rect 15102 14220 15108 14232
rect 15160 14220 15166 14272
rect 35802 14260 35808 14272
rect 35763 14232 35808 14260
rect 35802 14220 35808 14232
rect 35860 14220 35866 14272
rect 1104 14170 68816 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 68816 14170
rect 1104 14096 68816 14118
rect 30653 13991 30711 13997
rect 30653 13957 30665 13991
rect 30699 13988 30711 13991
rect 31938 13988 31944 14000
rect 30699 13960 31944 13988
rect 30699 13957 30711 13960
rect 30653 13951 30711 13957
rect 31938 13948 31944 13960
rect 31996 13948 32002 14000
rect 30742 13920 30748 13932
rect 30703 13892 30748 13920
rect 30742 13880 30748 13892
rect 30800 13880 30806 13932
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 12250 13852 12256 13864
rect 10735 13824 12256 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 31389 13855 31447 13861
rect 31389 13821 31401 13855
rect 31435 13852 31447 13855
rect 32122 13852 32128 13864
rect 31435 13824 32128 13852
rect 31435 13821 31447 13824
rect 31389 13815 31447 13821
rect 32122 13812 32128 13824
rect 32180 13812 32186 13864
rect 14918 13676 14924 13728
rect 14976 13716 14982 13728
rect 15013 13719 15071 13725
rect 15013 13716 15025 13719
rect 14976 13688 15025 13716
rect 14976 13676 14982 13688
rect 15013 13685 15025 13688
rect 15059 13685 15071 13719
rect 15013 13679 15071 13685
rect 1104 13626 68816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 68816 13626
rect 1104 13552 68816 13574
rect 36354 13444 36360 13456
rect 35636 13416 36360 13444
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 4120 13348 10425 13376
rect 4120 13336 4126 13348
rect 10413 13345 10425 13348
rect 10459 13345 10471 13379
rect 12250 13376 12256 13388
rect 12211 13348 12256 13376
rect 10413 13339 10471 13345
rect 12250 13336 12256 13348
rect 12308 13336 12314 13388
rect 14918 13376 14924 13388
rect 14879 13348 14924 13376
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 15102 13376 15108 13388
rect 15063 13348 15108 13376
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15470 13376 15476 13388
rect 15431 13348 15476 13376
rect 15470 13336 15476 13348
rect 15528 13336 15534 13388
rect 31938 13376 31944 13388
rect 31899 13348 31944 13376
rect 31938 13336 31944 13348
rect 31996 13336 32002 13388
rect 32122 13376 32128 13388
rect 32083 13348 32128 13376
rect 32122 13336 32128 13348
rect 32180 13336 32186 13388
rect 35636 13385 35664 13416
rect 36354 13404 36360 13416
rect 36412 13404 36418 13456
rect 35621 13379 35679 13385
rect 35621 13345 35633 13379
rect 35667 13345 35679 13379
rect 35802 13376 35808 13388
rect 35763 13348 35808 13376
rect 35621 13339 35679 13345
rect 35802 13336 35808 13348
rect 35860 13336 35866 13388
rect 36078 13376 36084 13388
rect 36039 13348 36084 13376
rect 36078 13336 36084 13348
rect 36136 13336 36142 13388
rect 11606 13200 11612 13252
rect 11664 13240 11670 13252
rect 12069 13243 12127 13249
rect 12069 13240 12081 13243
rect 11664 13212 12081 13240
rect 11664 13200 11670 13212
rect 12069 13209 12081 13212
rect 12115 13209 12127 13243
rect 30282 13240 30288 13252
rect 30243 13212 30288 13240
rect 12069 13203 12127 13209
rect 30282 13200 30288 13212
rect 30340 13200 30346 13252
rect 1104 13082 68816 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 68816 13082
rect 1104 13008 68816 13030
rect 11606 12968 11612 12980
rect 11567 12940 11612 12968
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 30282 12968 30288 12980
rect 12406 12940 30288 12968
rect 3326 12860 3332 12912
rect 3384 12900 3390 12912
rect 12406 12900 12434 12940
rect 30282 12928 30288 12940
rect 30340 12928 30346 12980
rect 3384 12872 12434 12900
rect 3384 12860 3390 12872
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12832 11759 12835
rect 11790 12832 11796 12844
rect 11747 12804 11796 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 9030 12628 9036 12640
rect 8991 12600 9036 12628
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 1104 12538 68816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 68816 12538
rect 1104 12464 68816 12486
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 8938 12220 8944 12232
rect 8343 12192 8944 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9674 12220 9680 12232
rect 9635 12192 9680 12220
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 40034 12180 40040 12232
rect 40092 12220 40098 12232
rect 40221 12223 40279 12229
rect 40221 12220 40233 12223
rect 40092 12192 40233 12220
rect 40092 12180 40098 12192
rect 40221 12189 40233 12192
rect 40267 12189 40279 12223
rect 41506 12220 41512 12232
rect 41467 12192 41512 12220
rect 40221 12183 40279 12189
rect 41506 12180 41512 12192
rect 41564 12180 41570 12232
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 9585 12087 9643 12093
rect 9585 12084 9597 12087
rect 9272 12056 9597 12084
rect 9272 12044 9278 12056
rect 9585 12053 9597 12056
rect 9631 12053 9643 12087
rect 9585 12047 9643 12053
rect 41601 12087 41659 12093
rect 41601 12053 41613 12087
rect 41647 12084 41659 12087
rect 41874 12084 41880 12096
rect 41647 12056 41880 12084
rect 41647 12053 41659 12056
rect 41601 12047 41659 12053
rect 41874 12044 41880 12056
rect 41932 12044 41938 12096
rect 1104 11994 68816 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 68816 11994
rect 1104 11920 68816 11942
rect 9214 11812 9220 11824
rect 9175 11784 9220 11812
rect 9214 11772 9220 11784
rect 9272 11772 9278 11824
rect 8386 11744 8392 11756
rect 8347 11716 8392 11744
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 9030 11744 9036 11756
rect 8991 11716 9036 11744
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 40034 11744 40040 11756
rect 39995 11716 40040 11744
rect 40034 11704 40040 11716
rect 40092 11704 40098 11756
rect 9766 11676 9772 11688
rect 9727 11648 9772 11676
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 40218 11676 40224 11688
rect 40179 11648 40224 11676
rect 40218 11636 40224 11648
rect 40276 11636 40282 11688
rect 41877 11679 41935 11685
rect 41877 11645 41889 11679
rect 41923 11676 41935 11679
rect 62114 11676 62120 11688
rect 41923 11648 62120 11676
rect 41923 11645 41935 11648
rect 41877 11639 41935 11645
rect 62114 11636 62120 11648
rect 62172 11636 62178 11688
rect 8481 11543 8539 11549
rect 8481 11509 8493 11543
rect 8527 11540 8539 11543
rect 9122 11540 9128 11552
rect 8527 11512 9128 11540
rect 8527 11509 8539 11512
rect 8481 11503 8539 11509
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 24394 11540 24400 11552
rect 24355 11512 24400 11540
rect 24394 11500 24400 11512
rect 24452 11500 24458 11552
rect 41690 11500 41696 11552
rect 41748 11540 41754 11552
rect 42429 11543 42487 11549
rect 42429 11540 42441 11543
rect 41748 11512 42441 11540
rect 41748 11500 41754 11512
rect 42429 11509 42441 11512
rect 42475 11509 42487 11543
rect 42429 11503 42487 11509
rect 1104 11450 68816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 68816 11450
rect 1104 11376 68816 11398
rect 40129 11339 40187 11345
rect 40129 11305 40141 11339
rect 40175 11336 40187 11339
rect 40218 11336 40224 11348
rect 40175 11308 40224 11336
rect 40175 11305 40187 11308
rect 40129 11299 40187 11305
rect 40218 11296 40224 11308
rect 40276 11296 40282 11348
rect 20714 11228 20720 11280
rect 20772 11268 20778 11280
rect 20772 11240 24900 11268
rect 20772 11228 20778 11240
rect 8938 11200 8944 11212
rect 8899 11172 8944 11200
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9122 11200 9128 11212
rect 9083 11172 9128 11200
rect 9122 11160 9128 11172
rect 9180 11160 9186 11212
rect 9858 11200 9864 11212
rect 9819 11172 9864 11200
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 24394 11200 24400 11212
rect 24355 11172 24400 11200
rect 24394 11160 24400 11172
rect 24452 11160 24458 11212
rect 24872 11209 24900 11240
rect 24857 11203 24915 11209
rect 24857 11169 24869 11203
rect 24903 11169 24915 11203
rect 41690 11200 41696 11212
rect 41651 11172 41696 11200
rect 24857 11163 24915 11169
rect 41690 11160 41696 11172
rect 41748 11160 41754 11212
rect 41874 11200 41880 11212
rect 41835 11172 41880 11200
rect 41874 11160 41880 11172
rect 41932 11160 41938 11212
rect 27522 11132 27528 11144
rect 27483 11104 27528 11132
rect 27522 11092 27528 11104
rect 27580 11092 27586 11144
rect 40037 11135 40095 11141
rect 40037 11101 40049 11135
rect 40083 11132 40095 11135
rect 40126 11132 40132 11144
rect 40083 11104 40132 11132
rect 40083 11101 40095 11104
rect 40037 11095 40095 11101
rect 40126 11092 40132 11104
rect 40184 11092 40190 11144
rect 24578 11064 24584 11076
rect 24539 11036 24584 11064
rect 24578 11024 24584 11036
rect 24636 11024 24642 11076
rect 43533 11067 43591 11073
rect 43533 11033 43545 11067
rect 43579 11064 43591 11067
rect 57238 11064 57244 11076
rect 43579 11036 57244 11064
rect 43579 11033 43591 11036
rect 43533 11027 43591 11033
rect 57238 11024 57244 11036
rect 57296 11024 57302 11076
rect 3418 10956 3424 11008
rect 3476 10996 3482 11008
rect 9766 10996 9772 11008
rect 3476 10968 9772 10996
rect 3476 10956 3482 10968
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 1104 10906 68816 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 68816 10906
rect 1104 10832 68816 10854
rect 24578 10752 24584 10804
rect 24636 10792 24642 10804
rect 24765 10795 24823 10801
rect 24765 10792 24777 10795
rect 24636 10764 24777 10792
rect 24636 10752 24642 10764
rect 24765 10761 24777 10764
rect 24811 10761 24823 10795
rect 24765 10755 24823 10761
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 9732 10628 10241 10656
rect 9732 10616 9738 10628
rect 10229 10625 10241 10628
rect 10275 10625 10287 10659
rect 24854 10656 24860 10668
rect 24815 10628 24860 10656
rect 10229 10619 10287 10625
rect 24854 10616 24860 10628
rect 24912 10616 24918 10668
rect 27522 10656 27528 10668
rect 27483 10628 27528 10656
rect 27522 10616 27528 10628
rect 27580 10616 27586 10668
rect 38194 10656 38200 10668
rect 38155 10628 38200 10656
rect 38194 10616 38200 10628
rect 38252 10616 38258 10668
rect 40126 10616 40132 10668
rect 40184 10656 40190 10668
rect 43993 10659 44051 10665
rect 43993 10656 44005 10659
rect 40184 10628 44005 10656
rect 40184 10616 40190 10628
rect 43993 10625 44005 10628
rect 44039 10625 44051 10659
rect 43993 10619 44051 10625
rect 62114 10616 62120 10668
rect 62172 10656 62178 10668
rect 66162 10656 66168 10668
rect 62172 10628 66168 10656
rect 62172 10616 62178 10628
rect 66162 10616 66168 10628
rect 66220 10616 66226 10668
rect 27709 10591 27767 10597
rect 27709 10557 27721 10591
rect 27755 10588 27767 10591
rect 27890 10588 27896 10600
rect 27755 10560 27896 10588
rect 27755 10557 27767 10560
rect 27709 10551 27767 10557
rect 27890 10548 27896 10560
rect 27948 10548 27954 10600
rect 29362 10588 29368 10600
rect 29323 10560 29368 10588
rect 29362 10548 29368 10560
rect 29420 10548 29426 10600
rect 9585 10455 9643 10461
rect 9585 10421 9597 10455
rect 9631 10452 9643 10455
rect 9766 10452 9772 10464
rect 9631 10424 9772 10452
rect 9631 10421 9643 10424
rect 9585 10415 9643 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10137 10455 10195 10461
rect 10137 10452 10149 10455
rect 10008 10424 10149 10452
rect 10008 10412 10014 10424
rect 10137 10421 10149 10424
rect 10183 10421 10195 10455
rect 38286 10452 38292 10464
rect 38247 10424 38292 10452
rect 10137 10415 10195 10421
rect 38286 10412 38292 10424
rect 38344 10412 38350 10464
rect 38838 10452 38844 10464
rect 38799 10424 38844 10452
rect 38838 10412 38844 10424
rect 38896 10412 38902 10464
rect 44082 10452 44088 10464
rect 44043 10424 44088 10452
rect 44082 10412 44088 10424
rect 44140 10412 44146 10464
rect 44821 10455 44879 10461
rect 44821 10421 44833 10455
rect 44867 10452 44879 10455
rect 45002 10452 45008 10464
rect 44867 10424 45008 10452
rect 44867 10421 44879 10424
rect 44821 10415 44879 10421
rect 45002 10412 45008 10424
rect 45060 10412 45066 10464
rect 1104 10362 68816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 68816 10362
rect 1104 10288 68816 10310
rect 27890 10248 27896 10260
rect 27851 10220 27896 10248
rect 27890 10208 27896 10220
rect 27948 10208 27954 10260
rect 44082 10140 44088 10192
rect 44140 10180 44146 10192
rect 44140 10152 45232 10180
rect 44140 10140 44146 10152
rect 9766 10112 9772 10124
rect 9727 10084 9772 10112
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 9950 10112 9956 10124
rect 9911 10084 9956 10112
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 10318 10112 10324 10124
rect 10279 10084 10324 10112
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 45002 10112 45008 10124
rect 44963 10084 45008 10112
rect 45002 10072 45008 10084
rect 45060 10072 45066 10124
rect 45204 10121 45232 10152
rect 45189 10115 45247 10121
rect 45189 10081 45201 10115
rect 45235 10081 45247 10115
rect 45189 10075 45247 10081
rect 24854 10004 24860 10056
rect 24912 10044 24918 10056
rect 27985 10047 28043 10053
rect 27985 10044 27997 10047
rect 24912 10016 27997 10044
rect 24912 10004 24918 10016
rect 27985 10013 27997 10016
rect 28031 10044 28043 10047
rect 38194 10044 38200 10056
rect 28031 10016 38200 10044
rect 28031 10013 28043 10016
rect 27985 10007 28043 10013
rect 38194 10004 38200 10016
rect 38252 10004 38258 10056
rect 46845 9979 46903 9985
rect 46845 9945 46857 9979
rect 46891 9976 46903 9979
rect 62758 9976 62764 9988
rect 46891 9948 62764 9976
rect 46891 9945 46903 9948
rect 46845 9939 46903 9945
rect 62758 9936 62764 9948
rect 62816 9936 62822 9988
rect 1104 9818 68816 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 68816 9818
rect 1104 9744 68816 9766
rect 3418 9596 3424 9648
rect 3476 9636 3482 9648
rect 9858 9636 9864 9648
rect 3476 9608 9864 9636
rect 3476 9596 3482 9608
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 38286 9636 38292 9648
rect 38247 9608 38292 9636
rect 38286 9596 38292 9608
rect 38344 9596 38350 9648
rect 38105 9503 38163 9509
rect 38105 9469 38117 9503
rect 38151 9469 38163 9503
rect 38654 9500 38660 9512
rect 38615 9472 38660 9500
rect 38105 9463 38163 9469
rect 38120 9432 38148 9463
rect 38654 9460 38660 9472
rect 38712 9460 38718 9512
rect 38838 9432 38844 9444
rect 38120 9404 38844 9432
rect 38838 9392 38844 9404
rect 38896 9392 38902 9444
rect 1104 9274 68816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 68816 9274
rect 1104 9200 68816 9222
rect 1104 8730 68816 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 68816 8730
rect 1104 8656 68816 8678
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 20714 8276 20720 8288
rect 3476 8248 20720 8276
rect 3476 8236 3482 8248
rect 20714 8236 20720 8248
rect 20772 8236 20778 8288
rect 47762 8236 47768 8288
rect 47820 8276 47826 8288
rect 47857 8279 47915 8285
rect 47857 8276 47869 8279
rect 47820 8248 47869 8276
rect 47820 8236 47826 8248
rect 47857 8245 47869 8248
rect 47903 8245 47915 8279
rect 47857 8239 47915 8245
rect 1104 8186 68816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 68816 8186
rect 1104 8112 68816 8134
rect 47762 7936 47768 7948
rect 47723 7908 47768 7936
rect 47762 7896 47768 7908
rect 47820 7896 47826 7948
rect 47118 7868 47124 7880
rect 47079 7840 47124 7868
rect 47118 7828 47124 7840
rect 47176 7828 47182 7880
rect 47213 7803 47271 7809
rect 47213 7769 47225 7803
rect 47259 7800 47271 7803
rect 47949 7803 48007 7809
rect 47949 7800 47961 7803
rect 47259 7772 47961 7800
rect 47259 7769 47271 7772
rect 47213 7763 47271 7769
rect 47949 7769 47961 7772
rect 47995 7769 48007 7803
rect 47949 7763 48007 7769
rect 49605 7803 49663 7809
rect 49605 7769 49617 7803
rect 49651 7800 49663 7803
rect 66162 7800 66168 7812
rect 49651 7772 66168 7800
rect 49651 7769 49663 7772
rect 49605 7763 49663 7769
rect 66162 7760 66168 7772
rect 66220 7760 66226 7812
rect 1104 7642 68816 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 68816 7642
rect 1104 7568 68816 7590
rect 1104 7098 68816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 68816 7098
rect 1104 7024 68816 7046
rect 43254 6808 43260 6860
rect 43312 6848 43318 6860
rect 47118 6848 47124 6860
rect 43312 6820 47124 6848
rect 43312 6808 43318 6820
rect 47118 6808 47124 6820
rect 47176 6808 47182 6860
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 11146 6780 11152 6792
rect 10919 6752 11152 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11333 6783 11391 6789
rect 11333 6749 11345 6783
rect 11379 6749 11391 6783
rect 11333 6743 11391 6749
rect 10778 6672 10784 6724
rect 10836 6712 10842 6724
rect 10962 6712 10968 6724
rect 10836 6684 10968 6712
rect 10836 6672 10842 6684
rect 10962 6672 10968 6684
rect 11020 6712 11026 6724
rect 11348 6712 11376 6743
rect 11514 6740 11520 6792
rect 11572 6780 11578 6792
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11572 6752 11989 6780
rect 11572 6740 11578 6752
rect 11977 6749 11989 6752
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 11020 6684 11376 6712
rect 11020 6672 11026 6684
rect 11425 6647 11483 6653
rect 11425 6613 11437 6647
rect 11471 6644 11483 6647
rect 11698 6644 11704 6656
rect 11471 6616 11704 6644
rect 11471 6613 11483 6616
rect 11425 6607 11483 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 1104 6554 68816 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 68816 6554
rect 1104 6480 68816 6502
rect 11698 6372 11704 6384
rect 11659 6344 11704 6372
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 10778 6304 10784 6316
rect 10739 6276 10784 6304
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 11514 6304 11520 6316
rect 11475 6276 11520 6304
rect 11514 6264 11520 6276
rect 11572 6264 11578 6316
rect 43254 6264 43260 6316
rect 43312 6304 43318 6316
rect 43349 6307 43407 6313
rect 43349 6304 43361 6307
rect 43312 6276 43361 6304
rect 43312 6264 43318 6276
rect 43349 6273 43361 6276
rect 43395 6273 43407 6307
rect 43349 6267 43407 6273
rect 12434 6236 12440 6248
rect 12395 6208 12440 6236
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 10873 6103 10931 6109
rect 10873 6069 10885 6103
rect 10919 6100 10931 6103
rect 11330 6100 11336 6112
rect 10919 6072 11336 6100
rect 10919 6069 10931 6072
rect 10873 6063 10931 6069
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 43441 6103 43499 6109
rect 43441 6069 43453 6103
rect 43487 6100 43499 6103
rect 43622 6100 43628 6112
rect 43487 6072 43628 6100
rect 43487 6069 43499 6072
rect 43441 6063 43499 6069
rect 43622 6060 43628 6072
rect 43680 6060 43686 6112
rect 1104 6010 68816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 68816 6010
rect 1104 5936 68816 5958
rect 9030 5788 9036 5840
rect 9088 5828 9094 5840
rect 9088 5800 11652 5828
rect 9088 5788 9094 5800
rect 11146 5760 11152 5772
rect 11107 5732 11152 5760
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 11330 5760 11336 5772
rect 11291 5732 11336 5760
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 11624 5769 11652 5800
rect 11609 5763 11667 5769
rect 11609 5729 11621 5763
rect 11655 5729 11667 5763
rect 11609 5723 11667 5729
rect 43438 5652 43444 5704
rect 43496 5692 43502 5704
rect 43533 5695 43591 5701
rect 43533 5692 43545 5695
rect 43496 5664 43545 5692
rect 43496 5652 43502 5664
rect 43533 5661 43545 5664
rect 43579 5661 43591 5695
rect 43533 5655 43591 5661
rect 1104 5466 68816 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 68816 5466
rect 1104 5392 68816 5414
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 12434 5352 12440 5364
rect 3476 5324 12440 5352
rect 3476 5312 3482 5324
rect 12434 5312 12440 5324
rect 12492 5312 12498 5364
rect 3142 5244 3148 5296
rect 3200 5284 3206 5296
rect 10318 5284 10324 5296
rect 3200 5256 10324 5284
rect 3200 5244 3206 5256
rect 10318 5244 10324 5256
rect 10376 5244 10382 5296
rect 43622 5284 43628 5296
rect 43583 5256 43628 5284
rect 43622 5244 43628 5256
rect 43680 5244 43686 5296
rect 43438 5216 43444 5228
rect 43399 5188 43444 5216
rect 43438 5176 43444 5188
rect 43496 5176 43502 5228
rect 45281 5151 45339 5157
rect 45281 5117 45293 5151
rect 45327 5148 45339 5151
rect 60642 5148 60648 5160
rect 45327 5120 60648 5148
rect 45327 5117 45339 5120
rect 45281 5111 45339 5117
rect 60642 5108 60648 5120
rect 60700 5108 60706 5160
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 13538 5012 13544 5024
rect 12483 4984 13544 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 1104 4922 68816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 68816 4922
rect 1104 4848 68816 4870
rect 28994 4700 29000 4752
rect 29052 4740 29058 4752
rect 29549 4743 29607 4749
rect 29549 4740 29561 4743
rect 29052 4712 29561 4740
rect 29052 4700 29058 4712
rect 29549 4709 29561 4712
rect 29595 4709 29607 4743
rect 29549 4703 29607 4709
rect 13538 4672 13544 4684
rect 13499 4644 13544 4672
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 28997 4607 29055 4613
rect 28997 4573 29009 4607
rect 29043 4604 29055 4607
rect 29546 4604 29552 4616
rect 29043 4576 29552 4604
rect 29043 4573 29055 4576
rect 28997 4567 29055 4573
rect 29546 4564 29552 4576
rect 29604 4564 29610 4616
rect 11606 4496 11612 4548
rect 11664 4536 11670 4548
rect 11701 4539 11759 4545
rect 11701 4536 11713 4539
rect 11664 4508 11713 4536
rect 11664 4496 11670 4508
rect 11701 4505 11713 4508
rect 11747 4505 11759 4539
rect 13354 4536 13360 4548
rect 13315 4508 13360 4536
rect 11701 4499 11759 4505
rect 13354 4496 13360 4508
rect 13412 4496 13418 4548
rect 1104 4378 68816 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 68816 4378
rect 1104 4304 68816 4326
rect 12529 4267 12587 4273
rect 12529 4233 12541 4267
rect 12575 4264 12587 4267
rect 13354 4264 13360 4276
rect 12575 4236 13360 4264
rect 12575 4233 12587 4236
rect 12529 4227 12587 4233
rect 13354 4224 13360 4236
rect 13412 4224 13418 4276
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12437 4131 12495 4137
rect 12437 4128 12449 4131
rect 11848 4100 12449 4128
rect 11848 4088 11854 4100
rect 12437 4097 12449 4100
rect 12483 4128 12495 4131
rect 28353 4131 28411 4137
rect 28353 4128 28365 4131
rect 12483 4100 28365 4128
rect 12483 4097 12495 4100
rect 12437 4091 12495 4097
rect 28353 4097 28365 4100
rect 28399 4128 28411 4131
rect 28810 4128 28816 4140
rect 28399 4100 28816 4128
rect 28399 4097 28411 4100
rect 28353 4091 28411 4097
rect 28810 4088 28816 4100
rect 28868 4088 28874 4140
rect 28994 4128 29000 4140
rect 28955 4100 29000 4128
rect 28994 4088 29000 4100
rect 29052 4088 29058 4140
rect 62758 4088 62764 4140
rect 62816 4128 62822 4140
rect 66162 4128 66168 4140
rect 62816 4100 66168 4128
rect 62816 4088 62822 4100
rect 66162 4088 66168 4100
rect 66220 4088 66226 4140
rect 29181 4063 29239 4069
rect 29181 4029 29193 4063
rect 29227 4029 29239 4063
rect 29638 4060 29644 4072
rect 29599 4032 29644 4060
rect 29181 4023 29239 4029
rect 28445 3995 28503 4001
rect 28445 3961 28457 3995
rect 28491 3992 28503 3995
rect 29196 3992 29224 4023
rect 29638 4020 29644 4032
rect 29696 4020 29702 4072
rect 28491 3964 29224 3992
rect 28491 3961 28503 3964
rect 28445 3955 28503 3961
rect 1104 3834 68816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 68816 3834
rect 1104 3760 68816 3782
rect 54570 3612 54576 3664
rect 54628 3652 54634 3664
rect 67634 3652 67640 3664
rect 54628 3624 67640 3652
rect 54628 3612 54634 3624
rect 67634 3612 67640 3624
rect 67692 3612 67698 3664
rect 24486 3544 24492 3596
rect 24544 3584 24550 3596
rect 29362 3584 29368 3596
rect 24544 3556 29368 3584
rect 24544 3544 24550 3556
rect 29362 3544 29368 3556
rect 29420 3544 29426 3596
rect 29546 3584 29552 3596
rect 29507 3556 29552 3584
rect 29546 3544 29552 3556
rect 29604 3544 29610 3596
rect 56042 3544 56048 3596
rect 56100 3584 56106 3596
rect 57330 3584 57336 3596
rect 56100 3556 57336 3584
rect 56100 3544 56106 3556
rect 57330 3544 57336 3556
rect 57388 3544 57394 3596
rect 57606 3544 57612 3596
rect 57664 3584 57670 3596
rect 58618 3584 58624 3596
rect 57664 3556 58624 3584
rect 57664 3544 57670 3556
rect 58618 3544 58624 3556
rect 58676 3544 58682 3596
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 14458 3516 14464 3528
rect 6512 3488 14464 3516
rect 6512 3476 6518 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 18046 3476 18052 3528
rect 18104 3516 18110 3528
rect 24118 3516 24124 3528
rect 18104 3488 24124 3516
rect 18104 3476 18110 3488
rect 24118 3476 24124 3488
rect 24176 3476 24182 3528
rect 28810 3516 28816 3528
rect 28771 3488 28816 3516
rect 28810 3476 28816 3488
rect 28868 3476 28874 3528
rect 37182 3476 37188 3528
rect 37240 3516 37246 3528
rect 68922 3516 68928 3528
rect 37240 3488 68928 3516
rect 37240 3476 37246 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 10318 3408 10324 3460
rect 10376 3448 10382 3460
rect 24670 3448 24676 3460
rect 10376 3420 24676 3448
rect 10376 3408 10382 3420
rect 24670 3408 24676 3420
rect 24728 3408 24734 3460
rect 28905 3451 28963 3457
rect 28905 3417 28917 3451
rect 28951 3448 28963 3451
rect 29733 3451 29791 3457
rect 29733 3448 29745 3451
rect 28951 3420 29745 3448
rect 28951 3417 28963 3420
rect 28905 3411 28963 3417
rect 29733 3417 29745 3420
rect 29779 3417 29791 3451
rect 29733 3411 29791 3417
rect 31389 3451 31447 3457
rect 31389 3417 31401 3451
rect 31435 3448 31447 3451
rect 65058 3448 65064 3460
rect 31435 3420 65064 3448
rect 31435 3417 31447 3420
rect 31389 3411 31447 3417
rect 65058 3408 65064 3420
rect 65116 3408 65122 3460
rect 57882 3340 57888 3392
rect 57940 3380 57946 3392
rect 59906 3380 59912 3392
rect 57940 3352 59912 3380
rect 57940 3340 57946 3352
rect 59906 3340 59912 3352
rect 59964 3340 59970 3392
rect 1104 3290 68816 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 68816 3290
rect 1104 3216 68816 3238
rect 60642 2796 60648 2848
rect 60700 2836 60706 2848
rect 63770 2836 63776 2848
rect 60700 2808 63776 2836
rect 60700 2796 60706 2808
rect 63770 2796 63776 2808
rect 63828 2796 63834 2848
rect 1104 2746 68816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 68816 2746
rect 1104 2672 68816 2694
rect 1104 2202 68816 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 68816 2202
rect 1104 2128 68816 2150
<< via1 >>
rect 19574 69606 19626 69658
rect 19638 69606 19690 69658
rect 19702 69606 19754 69658
rect 19766 69606 19818 69658
rect 19830 69606 19882 69658
rect 50294 69606 50346 69658
rect 50358 69606 50410 69658
rect 50422 69606 50474 69658
rect 50486 69606 50538 69658
rect 50550 69606 50602 69658
rect 62764 69164 62816 69216
rect 66076 69164 66128 69216
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 34934 69062 34986 69114
rect 34998 69062 35050 69114
rect 35062 69062 35114 69114
rect 35126 69062 35178 69114
rect 35190 69062 35242 69114
rect 65654 69062 65706 69114
rect 65718 69062 65770 69114
rect 65782 69062 65834 69114
rect 65846 69062 65898 69114
rect 65910 69062 65962 69114
rect 52828 68960 52880 69012
rect 56692 68960 56744 69012
rect 62028 68756 62080 68808
rect 65340 68756 65392 68808
rect 19574 68518 19626 68570
rect 19638 68518 19690 68570
rect 19702 68518 19754 68570
rect 19766 68518 19818 68570
rect 19830 68518 19882 68570
rect 50294 68518 50346 68570
rect 50358 68518 50410 68570
rect 50422 68518 50474 68570
rect 50486 68518 50538 68570
rect 50550 68518 50602 68570
rect 1952 68280 2004 68332
rect 15844 68280 15896 68332
rect 21272 68280 21324 68332
rect 35348 68280 35400 68332
rect 50620 68280 50672 68332
rect 66996 68280 67048 68332
rect 49424 68144 49476 68196
rect 54116 68144 54168 68196
rect 46848 68076 46900 68128
rect 51540 68076 51592 68128
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 34934 67974 34986 68026
rect 34998 67974 35050 68026
rect 35062 67974 35114 68026
rect 35126 67974 35178 68026
rect 35190 67974 35242 68026
rect 65654 67974 65706 68026
rect 65718 67974 65770 68026
rect 65782 67974 65834 68026
rect 65846 67974 65898 68026
rect 65910 67974 65962 68026
rect 48964 67872 49016 67924
rect 49884 67872 49936 67924
rect 19984 67736 20036 67788
rect 21272 67736 21324 67788
rect 19574 67430 19626 67482
rect 19638 67430 19690 67482
rect 19702 67430 19754 67482
rect 19766 67430 19818 67482
rect 19830 67430 19882 67482
rect 50294 67430 50346 67482
rect 50358 67430 50410 67482
rect 50422 67430 50474 67482
rect 50486 67430 50538 67482
rect 50550 67430 50602 67482
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 19574 66342 19626 66394
rect 19638 66342 19690 66394
rect 19702 66342 19754 66394
rect 19766 66342 19818 66394
rect 19830 66342 19882 66394
rect 50294 66342 50346 66394
rect 50358 66342 50410 66394
rect 50422 66342 50474 66394
rect 50486 66342 50538 66394
rect 50550 66342 50602 66394
rect 39212 66240 39264 66292
rect 65340 66240 65392 66292
rect 1400 66147 1452 66156
rect 1400 66113 1409 66147
rect 1409 66113 1443 66147
rect 1443 66113 1452 66147
rect 1400 66104 1452 66113
rect 1584 66079 1636 66088
rect 1584 66045 1593 66079
rect 1593 66045 1627 66079
rect 1627 66045 1636 66079
rect 1584 66036 1636 66045
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 19574 65254 19626 65306
rect 19638 65254 19690 65306
rect 19702 65254 19754 65306
rect 19766 65254 19818 65306
rect 19830 65254 19882 65306
rect 50294 65254 50346 65306
rect 50358 65254 50410 65306
rect 50422 65254 50474 65306
rect 50486 65254 50538 65306
rect 50550 65254 50602 65306
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 34934 64710 34986 64762
rect 34998 64710 35050 64762
rect 35062 64710 35114 64762
rect 35126 64710 35178 64762
rect 35190 64710 35242 64762
rect 65654 64710 65706 64762
rect 65718 64710 65770 64762
rect 65782 64710 65834 64762
rect 65846 64710 65898 64762
rect 65910 64710 65962 64762
rect 19432 64404 19484 64456
rect 19574 64166 19626 64218
rect 19638 64166 19690 64218
rect 19702 64166 19754 64218
rect 19766 64166 19818 64218
rect 19830 64166 19882 64218
rect 50294 64166 50346 64218
rect 50358 64166 50410 64218
rect 50422 64166 50474 64218
rect 50486 64166 50538 64218
rect 50550 64166 50602 64218
rect 21272 64039 21324 64048
rect 21272 64005 21281 64039
rect 21281 64005 21315 64039
rect 21315 64005 21324 64039
rect 21272 63996 21324 64005
rect 19432 63971 19484 63980
rect 19432 63937 19441 63971
rect 19441 63937 19475 63971
rect 19475 63937 19484 63971
rect 19432 63928 19484 63937
rect 20168 63860 20220 63912
rect 19340 63724 19392 63776
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 34934 63622 34986 63674
rect 34998 63622 35050 63674
rect 35062 63622 35114 63674
rect 35126 63622 35178 63674
rect 35190 63622 35242 63674
rect 65654 63622 65706 63674
rect 65718 63622 65770 63674
rect 65782 63622 65834 63674
rect 65846 63622 65898 63674
rect 65910 63622 65962 63674
rect 15844 63452 15896 63504
rect 19340 63427 19392 63436
rect 19340 63393 19349 63427
rect 19349 63393 19383 63427
rect 19383 63393 19392 63427
rect 19340 63384 19392 63393
rect 43352 63359 43404 63368
rect 43352 63325 43361 63359
rect 43361 63325 43395 63359
rect 43395 63325 43404 63359
rect 43352 63316 43404 63325
rect 43628 63316 43680 63368
rect 19432 63180 19484 63232
rect 43812 63180 43864 63232
rect 19574 63078 19626 63130
rect 19638 63078 19690 63130
rect 19702 63078 19754 63130
rect 19766 63078 19818 63130
rect 19830 63078 19882 63130
rect 50294 63078 50346 63130
rect 50358 63078 50410 63130
rect 50422 63078 50474 63130
rect 50486 63078 50538 63130
rect 50550 63078 50602 63130
rect 19432 62976 19484 63028
rect 20168 63019 20220 63028
rect 20168 62985 20177 63019
rect 20177 62985 20211 63019
rect 20211 62985 20220 63019
rect 20168 62976 20220 62985
rect 43812 62951 43864 62960
rect 43812 62917 43821 62951
rect 43821 62917 43855 62951
rect 43855 62917 43864 62951
rect 43812 62908 43864 62917
rect 43352 62840 43404 62892
rect 43628 62883 43680 62892
rect 43628 62849 43637 62883
rect 43637 62849 43671 62883
rect 43671 62849 43680 62883
rect 43628 62840 43680 62849
rect 48964 62772 49016 62824
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 34934 62534 34986 62586
rect 34998 62534 35050 62586
rect 35062 62534 35114 62586
rect 35126 62534 35178 62586
rect 35190 62534 35242 62586
rect 65654 62534 65706 62586
rect 65718 62534 65770 62586
rect 65782 62534 65834 62586
rect 65846 62534 65898 62586
rect 65910 62534 65962 62586
rect 32772 62271 32824 62280
rect 32772 62237 32781 62271
rect 32781 62237 32815 62271
rect 32815 62237 32824 62271
rect 32772 62228 32824 62237
rect 37280 62228 37332 62280
rect 5540 62160 5592 62212
rect 32588 62203 32640 62212
rect 32588 62169 32597 62203
rect 32597 62169 32631 62203
rect 32631 62169 32640 62203
rect 32588 62160 32640 62169
rect 19574 61990 19626 62042
rect 19638 61990 19690 62042
rect 19702 61990 19754 62042
rect 19766 61990 19818 62042
rect 19830 61990 19882 62042
rect 50294 61990 50346 62042
rect 50358 61990 50410 62042
rect 50422 61990 50474 62042
rect 50486 61990 50538 62042
rect 50550 61990 50602 62042
rect 32588 61888 32640 61940
rect 35624 61752 35676 61804
rect 54116 61820 54168 61872
rect 37280 61795 37332 61804
rect 37280 61761 37289 61795
rect 37289 61761 37323 61795
rect 37323 61761 37332 61795
rect 37280 61752 37332 61761
rect 32772 61684 32824 61736
rect 37372 61616 37424 61668
rect 45836 61548 45888 61600
rect 55312 61548 55364 61600
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 65654 61446 65706 61498
rect 65718 61446 65770 61498
rect 65782 61446 65834 61498
rect 65846 61446 65898 61498
rect 65910 61446 65962 61498
rect 45560 61276 45612 61328
rect 45836 61251 45888 61260
rect 45836 61217 45845 61251
rect 45845 61217 45879 61251
rect 45879 61217 45888 61251
rect 45836 61208 45888 61217
rect 55312 61251 55364 61260
rect 55312 61217 55321 61251
rect 55321 61217 55355 61251
rect 55355 61217 55364 61251
rect 55312 61208 55364 61217
rect 54116 61183 54168 61192
rect 54116 61149 54125 61183
rect 54125 61149 54159 61183
rect 54159 61149 54168 61183
rect 54116 61140 54168 61149
rect 46020 61115 46072 61124
rect 46020 61081 46029 61115
rect 46029 61081 46063 61115
rect 46063 61081 46072 61115
rect 46020 61072 46072 61081
rect 64880 61072 64932 61124
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 46020 60843 46072 60852
rect 46020 60809 46029 60843
rect 46029 60809 46063 60843
rect 46063 60809 46072 60843
rect 46020 60800 46072 60809
rect 3424 60732 3476 60784
rect 24860 60732 24912 60784
rect 45928 60707 45980 60716
rect 45928 60673 45937 60707
rect 45937 60673 45971 60707
rect 45971 60673 45980 60707
rect 45928 60664 45980 60673
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 65654 60358 65706 60410
rect 65718 60358 65770 60410
rect 65782 60358 65834 60410
rect 65846 60358 65898 60410
rect 65910 60358 65962 60410
rect 26976 60052 27028 60104
rect 35532 60052 35584 60104
rect 54852 60052 54904 60104
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 26240 59619 26292 59628
rect 26240 59585 26249 59619
rect 26249 59585 26283 59619
rect 26283 59585 26292 59619
rect 26976 59619 27028 59628
rect 26240 59576 26292 59585
rect 26976 59585 26985 59619
rect 26985 59585 27019 59619
rect 27019 59585 27028 59619
rect 26976 59576 27028 59585
rect 24860 59440 24912 59492
rect 62764 59644 62816 59696
rect 45928 59576 45980 59628
rect 54852 59619 54904 59628
rect 54852 59585 54861 59619
rect 54861 59585 54895 59619
rect 54895 59585 54904 59619
rect 54852 59576 54904 59585
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 65654 59270 65706 59322
rect 65718 59270 65770 59322
rect 65782 59270 65834 59322
rect 65846 59270 65898 59322
rect 65910 59270 65962 59322
rect 35532 59075 35584 59084
rect 35532 59041 35541 59075
rect 35541 59041 35575 59075
rect 35575 59041 35584 59075
rect 35532 59032 35584 59041
rect 37188 59075 37240 59084
rect 37188 59041 37197 59075
rect 37197 59041 37231 59075
rect 37231 59041 37240 59075
rect 37188 59032 37240 59041
rect 35716 58939 35768 58948
rect 35716 58905 35725 58939
rect 35725 58905 35759 58939
rect 35759 58905 35768 58939
rect 35716 58896 35768 58905
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 35716 58667 35768 58676
rect 35716 58633 35725 58667
rect 35725 58633 35759 58667
rect 35759 58633 35768 58667
rect 35716 58624 35768 58633
rect 66076 58556 66128 58608
rect 35440 58488 35492 58540
rect 40316 58488 40368 58540
rect 64512 58463 64564 58472
rect 38108 58352 38160 58404
rect 64512 58429 64521 58463
rect 64521 58429 64555 58463
rect 64555 58429 64564 58463
rect 64512 58420 64564 58429
rect 65524 58352 65576 58404
rect 37924 58284 37976 58336
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 65654 58182 65706 58234
rect 65718 58182 65770 58234
rect 65782 58182 65834 58234
rect 65846 58182 65898 58234
rect 65910 58182 65962 58234
rect 64512 58080 64564 58132
rect 65524 58080 65576 58132
rect 37924 57987 37976 57996
rect 37924 57953 37933 57987
rect 37933 57953 37967 57987
rect 37967 57953 37976 57987
rect 37924 57944 37976 57953
rect 40316 57944 40368 57996
rect 63684 57944 63736 57996
rect 34704 57919 34756 57928
rect 34704 57885 34713 57919
rect 34713 57885 34747 57919
rect 34747 57885 34756 57919
rect 34704 57876 34756 57885
rect 35348 57876 35400 57928
rect 38108 57919 38160 57928
rect 38108 57885 38117 57919
rect 38117 57885 38151 57919
rect 38151 57885 38160 57919
rect 63500 57919 63552 57928
rect 38108 57876 38160 57885
rect 63500 57885 63509 57919
rect 63509 57885 63543 57919
rect 63543 57885 63552 57919
rect 63500 57876 63552 57885
rect 64236 57740 64288 57792
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 34704 57468 34756 57520
rect 64236 57511 64288 57520
rect 64236 57477 64245 57511
rect 64245 57477 64279 57511
rect 64279 57477 64288 57511
rect 64236 57468 64288 57477
rect 66168 57468 66220 57520
rect 63500 57400 63552 57452
rect 34428 57375 34480 57384
rect 34428 57341 34437 57375
rect 34437 57341 34471 57375
rect 34471 57341 34480 57375
rect 34428 57332 34480 57341
rect 35808 57375 35860 57384
rect 35808 57341 35817 57375
rect 35817 57341 35851 57375
rect 35851 57341 35860 57375
rect 35808 57332 35860 57341
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 34428 56992 34480 57044
rect 35440 56788 35492 56840
rect 49240 56831 49292 56840
rect 49240 56797 49249 56831
rect 49249 56797 49283 56831
rect 49283 56797 49292 56831
rect 49240 56788 49292 56797
rect 63960 56788 64012 56840
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 63592 56448 63644 56500
rect 64420 56448 64472 56500
rect 49240 56355 49292 56364
rect 49240 56321 49249 56355
rect 49249 56321 49283 56355
rect 49283 56321 49292 56355
rect 49240 56312 49292 56321
rect 63960 56355 64012 56364
rect 63960 56321 63969 56355
rect 63969 56321 64003 56355
rect 64003 56321 64012 56355
rect 63960 56312 64012 56321
rect 2780 56244 2832 56296
rect 32956 56287 33008 56296
rect 32956 56253 32965 56287
rect 32965 56253 32999 56287
rect 32999 56253 33008 56287
rect 32956 56244 33008 56253
rect 33140 56287 33192 56296
rect 33140 56253 33149 56287
rect 33149 56253 33183 56287
rect 33183 56253 33192 56287
rect 33140 56244 33192 56253
rect 49240 56176 49292 56228
rect 64236 56244 64288 56296
rect 64420 56287 64472 56296
rect 64420 56253 64429 56287
rect 64429 56253 64463 56287
rect 64463 56253 64472 56287
rect 64420 56244 64472 56253
rect 66168 56176 66220 56228
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 32956 55947 33008 55956
rect 32956 55913 32965 55947
rect 32965 55913 32999 55947
rect 32999 55913 33008 55947
rect 32956 55904 33008 55913
rect 49240 55947 49292 55956
rect 49240 55913 49249 55947
rect 49249 55913 49283 55947
rect 49283 55913 49292 55947
rect 49240 55904 49292 55913
rect 64236 55947 64288 55956
rect 64236 55913 64245 55947
rect 64245 55913 64279 55947
rect 64279 55913 64288 55947
rect 64236 55904 64288 55913
rect 35348 55700 35400 55752
rect 35440 55700 35492 55752
rect 48688 55743 48740 55752
rect 48688 55709 48697 55743
rect 48697 55709 48731 55743
rect 48731 55709 48740 55743
rect 48688 55700 48740 55709
rect 63684 55743 63736 55752
rect 63684 55709 63693 55743
rect 63693 55709 63727 55743
rect 63727 55709 63736 55743
rect 63684 55700 63736 55709
rect 64696 55700 64748 55752
rect 64972 55700 65024 55752
rect 63592 55607 63644 55616
rect 63592 55573 63601 55607
rect 63601 55573 63635 55607
rect 63635 55573 63644 55607
rect 63592 55564 63644 55573
rect 65156 55564 65208 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 50620 55292 50672 55344
rect 65156 55335 65208 55344
rect 65156 55301 65165 55335
rect 65165 55301 65199 55335
rect 65199 55301 65208 55335
rect 65156 55292 65208 55301
rect 66812 55335 66864 55344
rect 66812 55301 66821 55335
rect 66821 55301 66855 55335
rect 66855 55301 66864 55335
rect 66812 55292 66864 55301
rect 3332 55224 3384 55276
rect 35348 55267 35400 55276
rect 35348 55233 35357 55267
rect 35357 55233 35391 55267
rect 35391 55233 35400 55267
rect 48688 55267 48740 55276
rect 35348 55224 35400 55233
rect 48688 55233 48697 55267
rect 48697 55233 48731 55267
rect 48731 55233 48740 55267
rect 48688 55224 48740 55233
rect 64972 55267 65024 55276
rect 64972 55233 64981 55267
rect 64981 55233 65015 55267
rect 65015 55233 65024 55267
rect 64972 55224 65024 55233
rect 34796 55156 34848 55208
rect 48872 55199 48924 55208
rect 48872 55165 48881 55199
rect 48881 55165 48915 55199
rect 48915 55165 48924 55199
rect 48872 55156 48924 55165
rect 63224 55020 63276 55072
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 33140 54816 33192 54868
rect 34796 54859 34848 54868
rect 34796 54825 34805 54859
rect 34805 54825 34839 54859
rect 34839 54825 34848 54859
rect 34796 54816 34848 54825
rect 48872 54816 48924 54868
rect 63224 54723 63276 54732
rect 63224 54689 63233 54723
rect 63233 54689 63267 54723
rect 63267 54689 63276 54723
rect 63224 54680 63276 54689
rect 63592 54680 63644 54732
rect 65064 54723 65116 54732
rect 65064 54689 65073 54723
rect 65073 54689 65107 54723
rect 65107 54689 65116 54723
rect 65064 54680 65116 54689
rect 38016 54612 38068 54664
rect 48596 54655 48648 54664
rect 48596 54621 48605 54655
rect 48605 54621 48639 54655
rect 48639 54621 48648 54655
rect 48596 54612 48648 54621
rect 40776 54544 40828 54596
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 40684 52844 40736 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 40132 52572 40184 52624
rect 40684 52547 40736 52556
rect 40684 52513 40693 52547
rect 40693 52513 40727 52547
rect 40727 52513 40736 52547
rect 40684 52504 40736 52513
rect 40868 52411 40920 52420
rect 40868 52377 40877 52411
rect 40877 52377 40911 52411
rect 40911 52377 40920 52411
rect 40868 52368 40920 52377
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 40868 52139 40920 52148
rect 40868 52105 40877 52139
rect 40877 52105 40911 52139
rect 40911 52105 40920 52139
rect 40868 52096 40920 52105
rect 40776 52003 40828 52012
rect 40776 51969 40785 52003
rect 40785 51969 40819 52003
rect 40819 51969 40828 52003
rect 40776 51960 40828 51969
rect 32312 51935 32364 51944
rect 32312 51901 32321 51935
rect 32321 51901 32355 51935
rect 32355 51901 32364 51935
rect 32312 51892 32364 51901
rect 31760 51824 31812 51876
rect 50988 51756 51040 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 32312 51552 32364 51604
rect 50988 51459 51040 51468
rect 50988 51425 50997 51459
rect 50997 51425 51031 51459
rect 51031 51425 51040 51459
rect 50988 51416 51040 51425
rect 52828 51459 52880 51468
rect 52828 51425 52837 51459
rect 52837 51425 52871 51459
rect 52871 51425 52880 51459
rect 52828 51416 52880 51425
rect 51172 51323 51224 51332
rect 51172 51289 51181 51323
rect 51181 51289 51215 51323
rect 51215 51289 51224 51323
rect 51172 51280 51224 51289
rect 37924 51212 37976 51264
rect 48596 51212 48648 51264
rect 48964 51212 49016 51264
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 51172 51008 51224 51060
rect 43444 50872 43496 50924
rect 24400 50668 24452 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 6920 50328 6972 50380
rect 24400 50303 24452 50312
rect 24400 50269 24409 50303
rect 24409 50269 24443 50303
rect 24443 50269 24452 50303
rect 24400 50260 24452 50269
rect 24860 50192 24912 50244
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 24860 49963 24912 49972
rect 24860 49929 24869 49963
rect 24869 49929 24903 49963
rect 24903 49929 24912 49963
rect 24860 49920 24912 49929
rect 35348 49784 35400 49836
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 54116 49172 54168 49224
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 51080 48696 51132 48748
rect 54116 48739 54168 48748
rect 54116 48705 54125 48739
rect 54125 48705 54159 48739
rect 54159 48705 54168 48739
rect 54116 48696 54168 48705
rect 65432 48628 65484 48680
rect 22652 48492 22704 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 22652 48195 22704 48204
rect 22652 48161 22661 48195
rect 22661 48161 22695 48195
rect 22695 48161 22704 48195
rect 22652 48152 22704 48161
rect 3700 48016 3752 48068
rect 21916 48016 21968 48068
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 21916 47787 21968 47796
rect 21916 47753 21925 47787
rect 21925 47753 21959 47787
rect 21959 47753 21968 47787
rect 21916 47744 21968 47753
rect 49424 47719 49476 47728
rect 49424 47685 49433 47719
rect 49433 47685 49467 47719
rect 49467 47685 49476 47719
rect 49424 47676 49476 47685
rect 22008 47651 22060 47660
rect 22008 47617 22017 47651
rect 22017 47617 22051 47651
rect 22051 47617 22060 47651
rect 22008 47608 22060 47617
rect 47768 47583 47820 47592
rect 47768 47549 47777 47583
rect 47777 47549 47811 47583
rect 47811 47549 47820 47583
rect 47768 47540 47820 47549
rect 61936 47447 61988 47456
rect 61936 47413 61945 47447
rect 61945 47413 61979 47447
rect 61979 47413 61988 47447
rect 61936 47404 61988 47413
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 47768 47200 47820 47252
rect 58072 47064 58124 47116
rect 66168 47132 66220 47184
rect 61936 47107 61988 47116
rect 61936 47073 61945 47107
rect 61945 47073 61979 47107
rect 61979 47073 61988 47107
rect 61936 47064 61988 47073
rect 64788 47064 64840 47116
rect 44916 46996 44968 47048
rect 40776 46928 40828 46980
rect 56508 46996 56560 47048
rect 62120 46971 62172 46980
rect 62120 46937 62129 46971
rect 62129 46937 62163 46971
rect 62163 46937 62172 46971
rect 62120 46928 62172 46937
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 62120 46656 62172 46708
rect 58072 46520 58124 46572
rect 60924 46520 60976 46572
rect 41420 46452 41472 46504
rect 42432 46452 42484 46504
rect 41972 46316 42024 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 35532 45908 35584 45960
rect 51080 46044 51132 46096
rect 41972 46019 42024 46028
rect 41972 45985 41981 46019
rect 41981 45985 42015 46019
rect 42015 45985 42024 46019
rect 41972 45976 42024 45985
rect 42432 46019 42484 46028
rect 42432 45985 42441 46019
rect 42441 45985 42475 46019
rect 42475 45985 42484 46019
rect 42432 45976 42484 45985
rect 61016 45951 61068 45960
rect 61016 45917 61025 45951
rect 61025 45917 61059 45951
rect 61059 45917 61068 45951
rect 61016 45908 61068 45917
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 61016 45500 61068 45552
rect 65984 45500 66036 45552
rect 60832 45407 60884 45416
rect 60832 45373 60841 45407
rect 60841 45373 60875 45407
rect 60875 45373 60884 45407
rect 60832 45364 60884 45373
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 60832 45024 60884 45076
rect 60556 44863 60608 44872
rect 60556 44829 60565 44863
rect 60565 44829 60599 44863
rect 60599 44829 60608 44863
rect 60556 44820 60608 44829
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 60280 43732 60332 43784
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 60280 43299 60332 43308
rect 60280 43265 60289 43299
rect 60289 43265 60323 43299
rect 60323 43265 60332 43299
rect 60280 43256 60332 43265
rect 60464 43231 60516 43240
rect 60464 43197 60473 43231
rect 60473 43197 60507 43231
rect 60507 43197 60516 43231
rect 60464 43188 60516 43197
rect 62028 43231 62080 43240
rect 62028 43197 62037 43231
rect 62037 43197 62071 43231
rect 62071 43197 62080 43231
rect 62028 43188 62080 43197
rect 16764 43052 16816 43104
rect 34704 43052 34756 43104
rect 45008 43052 45060 43104
rect 52736 43095 52788 43104
rect 52736 43061 52745 43095
rect 52745 43061 52779 43095
rect 52779 43061 52788 43095
rect 52736 43052 52788 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 60464 42848 60516 42900
rect 3700 42712 3752 42764
rect 45008 42755 45060 42764
rect 45008 42721 45017 42755
rect 45017 42721 45051 42755
rect 45051 42721 45060 42755
rect 45008 42712 45060 42721
rect 46848 42755 46900 42764
rect 46848 42721 46857 42755
rect 46857 42721 46891 42755
rect 46891 42721 46900 42755
rect 46848 42712 46900 42721
rect 52736 42712 52788 42764
rect 16764 42687 16816 42696
rect 16764 42653 16773 42687
rect 16773 42653 16807 42687
rect 16807 42653 16816 42687
rect 16764 42644 16816 42653
rect 34704 42687 34756 42696
rect 34704 42653 34713 42687
rect 34713 42653 34747 42687
rect 34747 42653 34756 42687
rect 34704 42644 34756 42653
rect 48964 42644 49016 42696
rect 59728 42644 59780 42696
rect 60556 42644 60608 42696
rect 16948 42619 17000 42628
rect 16948 42585 16957 42619
rect 16957 42585 16991 42619
rect 16991 42585 17000 42619
rect 16948 42576 17000 42585
rect 16580 42508 16632 42560
rect 34612 42576 34664 42628
rect 45008 42576 45060 42628
rect 66168 42576 66220 42628
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 16948 42347 17000 42356
rect 16948 42313 16957 42347
rect 16957 42313 16991 42347
rect 16991 42313 17000 42347
rect 16948 42304 17000 42313
rect 34612 42347 34664 42356
rect 34612 42313 34621 42347
rect 34621 42313 34655 42347
rect 34655 42313 34664 42347
rect 34612 42304 34664 42313
rect 45008 42347 45060 42356
rect 45008 42313 45017 42347
rect 45017 42313 45051 42347
rect 45051 42313 45060 42347
rect 45008 42304 45060 42313
rect 14464 42168 14516 42220
rect 32864 42168 32916 42220
rect 38200 42168 38252 42220
rect 44916 42211 44968 42220
rect 44916 42177 44925 42211
rect 44925 42177 44959 42211
rect 44959 42177 44968 42211
rect 44916 42168 44968 42177
rect 38844 42100 38896 42152
rect 57428 41964 57480 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 57428 41667 57480 41676
rect 57428 41633 57437 41667
rect 57437 41633 57471 41667
rect 57471 41633 57480 41667
rect 57428 41624 57480 41633
rect 59084 41667 59136 41676
rect 59084 41633 59093 41667
rect 59093 41633 59127 41667
rect 59127 41633 59136 41667
rect 59084 41624 59136 41633
rect 56784 41599 56836 41608
rect 56784 41565 56793 41599
rect 56793 41565 56827 41599
rect 56827 41565 56836 41599
rect 56784 41556 56836 41565
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 61384 40060 61436 40112
rect 66168 40060 66220 40112
rect 9772 39788 9824 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 3608 39312 3660 39364
rect 9772 39491 9824 39500
rect 9772 39457 9781 39491
rect 9781 39457 9815 39491
rect 9815 39457 9824 39491
rect 9772 39448 9824 39457
rect 32956 39380 33008 39432
rect 10416 39312 10468 39364
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 10416 39083 10468 39092
rect 10416 39049 10425 39083
rect 10425 39049 10459 39083
rect 10459 39049 10468 39083
rect 10416 39040 10468 39049
rect 10508 38947 10560 38956
rect 10508 38913 10517 38947
rect 10517 38913 10551 38947
rect 10551 38913 10560 38947
rect 10508 38904 10560 38913
rect 32956 38947 33008 38956
rect 32956 38913 32965 38947
rect 32965 38913 32999 38947
rect 32999 38913 33008 38947
rect 32956 38904 33008 38913
rect 64696 38947 64748 38956
rect 64696 38913 64705 38947
rect 64705 38913 64739 38947
rect 64739 38913 64748 38947
rect 64696 38904 64748 38913
rect 33140 38879 33192 38888
rect 33140 38845 33149 38879
rect 33149 38845 33183 38879
rect 33183 38845 33192 38879
rect 33140 38836 33192 38845
rect 65156 38836 65208 38888
rect 65340 38879 65392 38888
rect 65340 38845 65349 38879
rect 65349 38845 65383 38879
rect 65383 38845 65392 38879
rect 65340 38836 65392 38845
rect 67180 38879 67232 38888
rect 67180 38845 67189 38879
rect 67189 38845 67223 38879
rect 67223 38845 67232 38879
rect 67180 38836 67232 38845
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 33140 38496 33192 38548
rect 65340 38496 65392 38548
rect 32864 38335 32916 38344
rect 32864 38301 32873 38335
rect 32873 38301 32907 38335
rect 32907 38301 32916 38335
rect 32864 38292 32916 38301
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 37372 37655 37424 37664
rect 37372 37621 37381 37655
rect 37381 37621 37415 37655
rect 37415 37621 37424 37655
rect 37372 37612 37424 37621
rect 61660 37655 61712 37664
rect 61660 37621 61669 37655
rect 61669 37621 61703 37655
rect 61703 37621 61712 37655
rect 61660 37612 61712 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 37372 37315 37424 37324
rect 37372 37281 37381 37315
rect 37381 37281 37415 37315
rect 37415 37281 37424 37315
rect 37372 37272 37424 37281
rect 61660 37315 61712 37324
rect 61660 37281 61669 37315
rect 61669 37281 61703 37315
rect 61703 37281 61712 37315
rect 61660 37272 61712 37281
rect 66168 37272 66220 37324
rect 39212 37247 39264 37256
rect 32404 37179 32456 37188
rect 32404 37145 32413 37179
rect 32413 37145 32447 37179
rect 32447 37145 32456 37179
rect 32404 37136 32456 37145
rect 39212 37213 39221 37247
rect 39221 37213 39255 37247
rect 39255 37213 39264 37247
rect 39212 37204 39264 37213
rect 60924 37204 60976 37256
rect 61292 37204 61344 37256
rect 36544 37136 36596 37188
rect 36636 37136 36688 37188
rect 32496 37111 32548 37120
rect 32496 37077 32505 37111
rect 32505 37077 32539 37111
rect 32539 37077 32548 37111
rect 32496 37068 32548 37077
rect 37372 37068 37424 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 36636 36907 36688 36916
rect 36636 36873 36645 36907
rect 36645 36873 36679 36907
rect 36679 36873 36688 36907
rect 36636 36864 36688 36873
rect 1584 36796 1636 36848
rect 32404 36796 32456 36848
rect 32496 36796 32548 36848
rect 35624 36796 35676 36848
rect 34152 36728 34204 36780
rect 36084 36728 36136 36780
rect 37648 36796 37700 36848
rect 37924 36839 37976 36848
rect 37924 36805 37933 36839
rect 37933 36805 37967 36839
rect 37967 36805 37976 36839
rect 37924 36796 37976 36805
rect 38016 36796 38068 36848
rect 40316 36839 40368 36848
rect 40316 36805 40325 36839
rect 40325 36805 40359 36839
rect 40359 36805 40368 36839
rect 40316 36796 40368 36805
rect 37372 36771 37424 36780
rect 37372 36737 37381 36771
rect 37381 36737 37415 36771
rect 37415 36737 37424 36771
rect 37372 36728 37424 36737
rect 38660 36728 38712 36780
rect 64696 36728 64748 36780
rect 14188 36660 14240 36712
rect 13820 36592 13872 36644
rect 34704 36660 34756 36712
rect 35440 36660 35492 36712
rect 34428 36524 34480 36576
rect 64880 36567 64932 36576
rect 64880 36533 64889 36567
rect 64889 36533 64923 36567
rect 64923 36533 64932 36567
rect 64880 36524 64932 36533
rect 65524 36524 65576 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 14188 36363 14240 36372
rect 14188 36329 14197 36363
rect 14197 36329 14231 36363
rect 14231 36329 14240 36363
rect 14188 36320 14240 36329
rect 32956 36320 33008 36372
rect 43352 36320 43404 36372
rect 25320 36252 25372 36304
rect 64880 36252 64932 36304
rect 43444 36184 43496 36236
rect 65524 36184 65576 36236
rect 6368 36159 6420 36168
rect 6368 36125 6377 36159
rect 6377 36125 6411 36159
rect 6411 36125 6420 36159
rect 6368 36116 6420 36125
rect 14280 36159 14332 36168
rect 14280 36125 14289 36159
rect 14289 36125 14323 36159
rect 14323 36125 14332 36159
rect 14280 36116 14332 36125
rect 32496 36116 32548 36168
rect 33784 36159 33836 36168
rect 33784 36125 33793 36159
rect 33793 36125 33827 36159
rect 33827 36125 33836 36159
rect 33784 36116 33836 36125
rect 34152 36116 34204 36168
rect 36084 36159 36136 36168
rect 36084 36125 36093 36159
rect 36093 36125 36127 36159
rect 36127 36125 36136 36159
rect 36084 36116 36136 36125
rect 36544 36159 36596 36168
rect 36544 36125 36553 36159
rect 36553 36125 36587 36159
rect 36587 36125 36596 36159
rect 36544 36116 36596 36125
rect 37372 36116 37424 36168
rect 45192 36116 45244 36168
rect 32772 36048 32824 36100
rect 32956 36091 33008 36100
rect 32956 36057 32965 36091
rect 32965 36057 32999 36091
rect 32999 36057 33008 36091
rect 32956 36048 33008 36057
rect 26240 35980 26292 36032
rect 35440 35980 35492 36032
rect 35900 35980 35952 36032
rect 67456 36091 67508 36100
rect 67456 36057 67465 36091
rect 67465 36057 67499 36091
rect 67499 36057 67508 36091
rect 67456 36048 67508 36057
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 40684 35708 40736 35760
rect 61384 35708 61436 35760
rect 6368 35683 6420 35692
rect 6368 35649 6377 35683
rect 6377 35649 6411 35683
rect 6411 35649 6420 35683
rect 6368 35640 6420 35649
rect 32496 35640 32548 35692
rect 35900 35683 35952 35692
rect 35900 35649 35909 35683
rect 35909 35649 35943 35683
rect 35943 35649 35952 35683
rect 35900 35640 35952 35649
rect 41420 35640 41472 35692
rect 45192 35683 45244 35692
rect 45192 35649 45201 35683
rect 45201 35649 45235 35683
rect 45235 35649 45244 35683
rect 45192 35640 45244 35649
rect 6552 35615 6604 35624
rect 6552 35581 6561 35615
rect 6561 35581 6595 35615
rect 6595 35581 6604 35615
rect 6552 35572 6604 35581
rect 4068 35504 4120 35556
rect 14280 35572 14332 35624
rect 34612 35572 34664 35624
rect 35348 35615 35400 35624
rect 35348 35581 35357 35615
rect 35357 35581 35391 35615
rect 35391 35581 35400 35615
rect 35348 35572 35400 35581
rect 61292 35572 61344 35624
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 6552 35232 6604 35284
rect 6552 35071 6604 35080
rect 6552 35037 6561 35071
rect 6561 35037 6595 35071
rect 6595 35037 6604 35071
rect 6552 35028 6604 35037
rect 14280 35028 14332 35080
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 34796 34552 34848 34604
rect 35348 34552 35400 34604
rect 35900 34595 35952 34604
rect 35900 34561 35909 34595
rect 35909 34561 35943 34595
rect 35943 34561 35952 34595
rect 37372 34595 37424 34604
rect 35900 34552 35952 34561
rect 37372 34561 37381 34595
rect 37381 34561 37415 34595
rect 37415 34561 37424 34595
rect 37372 34552 37424 34561
rect 10508 34484 10560 34536
rect 10968 34484 11020 34536
rect 43260 34552 43312 34604
rect 38200 34484 38252 34536
rect 22008 34416 22060 34468
rect 25320 34416 25372 34468
rect 24860 34391 24912 34400
rect 24860 34357 24869 34391
rect 24869 34357 24903 34391
rect 24903 34357 24912 34391
rect 24860 34348 24912 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 3424 33872 3476 33924
rect 24860 34051 24912 34060
rect 24860 34017 24869 34051
rect 24869 34017 24903 34051
rect 24903 34017 24912 34051
rect 24860 34008 24912 34017
rect 35532 34008 35584 34060
rect 36452 34008 36504 34060
rect 41420 34008 41472 34060
rect 35900 33940 35952 33992
rect 37372 33940 37424 33992
rect 49148 33940 49200 33992
rect 55496 33940 55548 33992
rect 25228 33872 25280 33924
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 25228 33643 25280 33652
rect 25228 33609 25237 33643
rect 25237 33609 25271 33643
rect 25271 33609 25280 33643
rect 25228 33600 25280 33609
rect 25320 33507 25372 33516
rect 25320 33473 25329 33507
rect 25329 33473 25363 33507
rect 25363 33473 25372 33507
rect 25320 33464 25372 33473
rect 43352 33532 43404 33584
rect 42432 33439 42484 33448
rect 42432 33405 42441 33439
rect 42441 33405 42475 33439
rect 42475 33405 42484 33439
rect 42432 33396 42484 33405
rect 66076 33532 66128 33584
rect 49148 33507 49200 33516
rect 49148 33473 49157 33507
rect 49157 33473 49191 33507
rect 49191 33473 49200 33507
rect 49148 33464 49200 33473
rect 55496 33507 55548 33516
rect 55496 33473 55505 33507
rect 55505 33473 55539 33507
rect 55539 33473 55548 33507
rect 55496 33464 55548 33473
rect 49332 33439 49384 33448
rect 49332 33405 49341 33439
rect 49341 33405 49375 33439
rect 49375 33405 49384 33439
rect 49332 33396 49384 33405
rect 55680 33439 55732 33448
rect 55680 33405 55689 33439
rect 55689 33405 55723 33439
rect 55723 33405 55732 33439
rect 55680 33396 55732 33405
rect 57336 33439 57388 33448
rect 57336 33405 57345 33439
rect 57345 33405 57379 33439
rect 57379 33405 57388 33439
rect 57336 33396 57388 33405
rect 66168 33328 66220 33380
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 42432 33056 42484 33108
rect 49332 33056 49384 33108
rect 55680 33056 55732 33108
rect 40316 32852 40368 32904
rect 49056 32895 49108 32904
rect 49056 32861 49065 32895
rect 49065 32861 49099 32895
rect 49099 32861 49108 32895
rect 49056 32852 49108 32861
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 43444 32376 43496 32428
rect 49056 32512 49108 32564
rect 44548 32351 44600 32360
rect 44548 32317 44557 32351
rect 44557 32317 44591 32351
rect 44591 32317 44600 32351
rect 44548 32308 44600 32317
rect 44180 32240 44232 32292
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 44548 31968 44600 32020
rect 5448 31807 5500 31816
rect 5448 31773 5457 31807
rect 5457 31773 5491 31807
rect 5491 31773 5500 31807
rect 5448 31764 5500 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 6552 31331 6604 31340
rect 6552 31297 6561 31331
rect 6561 31297 6595 31331
rect 6595 31297 6604 31331
rect 6552 31288 6604 31297
rect 34428 31288 34480 31340
rect 38568 31288 38620 31340
rect 38844 31263 38896 31272
rect 38844 31229 38853 31263
rect 38853 31229 38887 31263
rect 38887 31229 38896 31263
rect 38844 31220 38896 31229
rect 56784 31220 56836 31272
rect 58164 31220 58216 31272
rect 5632 31084 5684 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 2964 30812 3016 30864
rect 5448 30787 5500 30796
rect 5448 30753 5457 30787
rect 5457 30753 5491 30787
rect 5491 30753 5500 30787
rect 5448 30744 5500 30753
rect 5632 30787 5684 30796
rect 5632 30753 5641 30787
rect 5641 30753 5675 30787
rect 5675 30753 5684 30787
rect 5632 30744 5684 30753
rect 32864 30787 32916 30796
rect 32864 30753 32873 30787
rect 32873 30753 32907 30787
rect 32907 30753 32916 30787
rect 32864 30744 32916 30753
rect 7748 30676 7800 30728
rect 19432 30676 19484 30728
rect 27988 30676 28040 30728
rect 33600 30676 33652 30728
rect 34428 30676 34480 30728
rect 59728 30719 59780 30728
rect 59728 30685 59737 30719
rect 59737 30685 59771 30719
rect 59771 30685 59780 30719
rect 59728 30676 59780 30685
rect 60464 30719 60516 30728
rect 60464 30685 60473 30719
rect 60473 30685 60507 30719
rect 60507 30685 60516 30719
rect 60464 30676 60516 30685
rect 66168 30608 66220 30660
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 7748 30243 7800 30252
rect 7748 30209 7757 30243
rect 7757 30209 7791 30243
rect 7791 30209 7800 30243
rect 7748 30200 7800 30209
rect 19432 30243 19484 30252
rect 19432 30209 19441 30243
rect 19441 30209 19475 30243
rect 19475 30209 19484 30243
rect 19432 30200 19484 30209
rect 27804 30200 27856 30252
rect 27988 30243 28040 30252
rect 27988 30209 27997 30243
rect 27997 30209 28031 30243
rect 28031 30209 28040 30243
rect 27988 30200 28040 30209
rect 60464 30200 60516 30252
rect 8300 30132 8352 30184
rect 3608 30064 3660 30116
rect 19984 30132 20036 30184
rect 19340 30064 19392 30116
rect 28356 30132 28408 30184
rect 26240 30064 26292 30116
rect 25504 30039 25556 30048
rect 25504 30005 25513 30039
rect 25513 30005 25547 30039
rect 25547 30005 25556 30039
rect 25504 29996 25556 30005
rect 25688 29996 25740 30048
rect 27528 30039 27580 30048
rect 27528 30005 27537 30039
rect 27537 30005 27571 30039
rect 27571 30005 27580 30039
rect 27528 29996 27580 30005
rect 51080 29996 51132 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 8300 29835 8352 29844
rect 8300 29801 8309 29835
rect 8309 29801 8343 29835
rect 8343 29801 8352 29835
rect 8300 29792 8352 29801
rect 19984 29835 20036 29844
rect 19984 29801 19993 29835
rect 19993 29801 20027 29835
rect 20027 29801 20036 29835
rect 19984 29792 20036 29801
rect 23480 29792 23532 29844
rect 28356 29835 28408 29844
rect 25504 29699 25556 29708
rect 25504 29665 25513 29699
rect 25513 29665 25547 29699
rect 25547 29665 25556 29699
rect 25504 29656 25556 29665
rect 25688 29699 25740 29708
rect 25688 29665 25697 29699
rect 25697 29665 25731 29699
rect 25731 29665 25740 29699
rect 25688 29656 25740 29665
rect 28356 29801 28365 29835
rect 28365 29801 28399 29835
rect 28399 29801 28408 29835
rect 28356 29792 28408 29801
rect 26056 29724 26108 29776
rect 32772 29724 32824 29776
rect 27804 29656 27856 29708
rect 8392 29631 8444 29640
rect 8392 29597 8401 29631
rect 8401 29597 8435 29631
rect 8435 29597 8444 29631
rect 8392 29588 8444 29597
rect 37648 29656 37700 29708
rect 35624 29588 35676 29640
rect 50988 29588 51040 29640
rect 26056 29520 26108 29572
rect 51724 29563 51776 29572
rect 51724 29529 51733 29563
rect 51733 29529 51767 29563
rect 51767 29529 51776 29563
rect 51724 29520 51776 29529
rect 53380 29563 53432 29572
rect 53380 29529 53389 29563
rect 53389 29529 53423 29563
rect 53423 29529 53432 29563
rect 53380 29520 53432 29529
rect 51264 29452 51316 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 35440 29248 35492 29300
rect 17960 29180 18012 29232
rect 38660 29248 38712 29300
rect 59728 29248 59780 29300
rect 27528 29155 27580 29164
rect 27528 29121 27537 29155
rect 27537 29121 27571 29155
rect 27571 29121 27580 29155
rect 27528 29112 27580 29121
rect 33784 29112 33836 29164
rect 27712 29087 27764 29096
rect 27712 29053 27721 29087
rect 27721 29053 27755 29087
rect 27755 29053 27764 29087
rect 27712 29044 27764 29053
rect 30748 29044 30800 29096
rect 38568 29112 38620 29164
rect 51724 29180 51776 29232
rect 28080 28976 28132 29028
rect 61660 29044 61712 29096
rect 38660 28976 38712 29028
rect 50988 29019 51040 29028
rect 50988 28985 50997 29019
rect 50997 28985 51031 29019
rect 51031 28985 51040 29019
rect 50988 28976 51040 28985
rect 3424 28908 3476 28960
rect 23480 28908 23532 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 27712 28704 27764 28756
rect 51080 28611 51132 28620
rect 51080 28577 51089 28611
rect 51089 28577 51123 28611
rect 51123 28577 51132 28611
rect 51080 28568 51132 28577
rect 51264 28611 51316 28620
rect 51264 28577 51273 28611
rect 51273 28577 51307 28611
rect 51307 28577 51316 28611
rect 51264 28568 51316 28577
rect 30748 28500 30800 28552
rect 33600 28543 33652 28552
rect 33600 28509 33609 28543
rect 33609 28509 33643 28543
rect 33643 28509 33652 28543
rect 33600 28500 33652 28509
rect 60648 28500 60700 28552
rect 8392 28432 8444 28484
rect 9128 28432 9180 28484
rect 40132 28432 40184 28484
rect 52920 28475 52972 28484
rect 52920 28441 52929 28475
rect 52929 28441 52963 28475
rect 52963 28441 52972 28475
rect 52920 28432 52972 28441
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 60648 28067 60700 28076
rect 60648 28033 60657 28067
rect 60657 28033 60691 28067
rect 60691 28033 60700 28067
rect 60648 28024 60700 28033
rect 50528 27999 50580 28008
rect 50528 27965 50537 27999
rect 50537 27965 50571 27999
rect 50571 27965 50580 27999
rect 50528 27956 50580 27965
rect 60832 27999 60884 28008
rect 60832 27965 60841 27999
rect 60841 27965 60875 27999
rect 60875 27965 60884 27999
rect 60832 27956 60884 27965
rect 64972 27956 65024 28008
rect 66168 27888 66220 27940
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 50528 27659 50580 27668
rect 50528 27625 50537 27659
rect 50537 27625 50571 27659
rect 50571 27625 50580 27659
rect 50528 27616 50580 27625
rect 60832 27616 60884 27668
rect 34704 27548 34756 27600
rect 35348 27548 35400 27600
rect 35532 27412 35584 27464
rect 61292 27455 61344 27464
rect 61292 27421 61301 27455
rect 61301 27421 61335 27455
rect 61335 27421 61344 27455
rect 61292 27412 61344 27421
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 33784 26911 33836 26920
rect 33784 26877 33793 26911
rect 33793 26877 33827 26911
rect 33827 26877 33836 26911
rect 33784 26868 33836 26877
rect 34796 26868 34848 26920
rect 6920 26800 6972 26852
rect 55772 26732 55824 26784
rect 58072 26732 58124 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 33784 26571 33836 26580
rect 33784 26537 33793 26571
rect 33793 26537 33827 26571
rect 33827 26537 33836 26571
rect 33784 26528 33836 26537
rect 34796 26571 34848 26580
rect 34796 26537 34805 26571
rect 34805 26537 34839 26571
rect 34839 26537 34848 26571
rect 34796 26528 34848 26537
rect 55772 26435 55824 26444
rect 55772 26401 55781 26435
rect 55781 26401 55815 26435
rect 55815 26401 55824 26435
rect 55772 26392 55824 26401
rect 58072 26435 58124 26444
rect 58072 26401 58081 26435
rect 58081 26401 58115 26435
rect 58115 26401 58124 26435
rect 58072 26392 58124 26401
rect 26884 26324 26936 26376
rect 35348 26324 35400 26376
rect 66168 26324 66220 26376
rect 55956 26299 56008 26308
rect 55956 26265 55965 26299
rect 55965 26265 55999 26299
rect 55999 26265 56008 26299
rect 55956 26256 56008 26265
rect 57612 26299 57664 26308
rect 57612 26265 57621 26299
rect 57621 26265 57655 26299
rect 57655 26265 57664 26299
rect 57612 26256 57664 26265
rect 58256 26299 58308 26308
rect 58256 26265 58265 26299
rect 58265 26265 58299 26299
rect 58299 26265 58308 26299
rect 58256 26256 58308 26265
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 55956 25984 56008 26036
rect 58256 26027 58308 26036
rect 58256 25993 58265 26027
rect 58265 25993 58299 26027
rect 58299 25993 58308 26027
rect 58256 25984 58308 25993
rect 27160 25891 27212 25900
rect 27160 25857 27169 25891
rect 27169 25857 27203 25891
rect 27203 25857 27212 25891
rect 27160 25848 27212 25857
rect 56508 25891 56560 25900
rect 56508 25857 56517 25891
rect 56517 25857 56551 25891
rect 56551 25857 56560 25891
rect 56508 25848 56560 25857
rect 58164 25891 58216 25900
rect 58164 25857 58173 25891
rect 58173 25857 58207 25891
rect 58207 25857 58216 25891
rect 58164 25848 58216 25857
rect 27528 25644 27580 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 26884 25372 26936 25424
rect 27528 25347 27580 25356
rect 27528 25313 27537 25347
rect 27537 25313 27571 25347
rect 27571 25313 27580 25347
rect 27528 25304 27580 25313
rect 32128 25304 32180 25356
rect 12348 25279 12400 25288
rect 12348 25245 12357 25279
rect 12357 25245 12391 25279
rect 12391 25245 12400 25279
rect 12348 25236 12400 25245
rect 28172 25279 28224 25288
rect 28172 25245 28181 25279
rect 28181 25245 28215 25279
rect 28215 25245 28224 25279
rect 28172 25236 28224 25245
rect 35716 25236 35768 25288
rect 3148 25168 3200 25220
rect 32312 25100 32364 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 27160 24896 27212 24948
rect 33692 24896 33744 24948
rect 32312 24871 32364 24880
rect 32312 24837 32321 24871
rect 32321 24837 32355 24871
rect 32355 24837 32364 24871
rect 32312 24828 32364 24837
rect 12348 24803 12400 24812
rect 12348 24769 12357 24803
rect 12357 24769 12391 24803
rect 12391 24769 12400 24803
rect 12348 24760 12400 24769
rect 27988 24760 28040 24812
rect 28172 24803 28224 24812
rect 28172 24769 28181 24803
rect 28181 24769 28215 24803
rect 28215 24769 28224 24803
rect 28172 24760 28224 24769
rect 32128 24803 32180 24812
rect 32128 24769 32137 24803
rect 32137 24769 32171 24803
rect 32171 24769 32180 24803
rect 32128 24760 32180 24769
rect 12992 24692 13044 24744
rect 3424 24624 3476 24676
rect 28540 24692 28592 24744
rect 3608 24556 3660 24608
rect 31760 24624 31812 24676
rect 23020 24599 23072 24608
rect 23020 24565 23029 24599
rect 23029 24565 23063 24599
rect 23063 24565 23072 24599
rect 23020 24556 23072 24565
rect 23204 24556 23256 24608
rect 27988 24556 28040 24608
rect 35440 24556 35492 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 12992 24395 13044 24404
rect 12992 24361 13001 24395
rect 13001 24361 13035 24395
rect 13035 24361 13044 24395
rect 12992 24352 13044 24361
rect 28540 24395 28592 24404
rect 28540 24361 28549 24395
rect 28549 24361 28583 24395
rect 28583 24361 28592 24395
rect 28540 24352 28592 24361
rect 14280 24148 14332 24200
rect 14464 24148 14516 24200
rect 34796 24148 34848 24200
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 23204 23783 23256 23792
rect 23204 23749 23213 23783
rect 23213 23749 23247 23783
rect 23247 23749 23256 23783
rect 23204 23740 23256 23749
rect 23020 23715 23072 23724
rect 23020 23681 23029 23715
rect 23029 23681 23063 23715
rect 23063 23681 23072 23715
rect 23020 23672 23072 23681
rect 24676 23647 24728 23656
rect 24676 23613 24685 23647
rect 24685 23613 24719 23647
rect 24719 23613 24728 23647
rect 24676 23604 24728 23613
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 35348 22584 35400 22636
rect 52184 22516 52236 22568
rect 54576 22559 54628 22568
rect 54576 22525 54585 22559
rect 54585 22525 54619 22559
rect 54619 22525 54628 22559
rect 54576 22516 54628 22525
rect 7564 22380 7616 22432
rect 9312 22423 9364 22432
rect 9312 22389 9321 22423
rect 9321 22389 9355 22423
rect 9355 22389 9364 22423
rect 9312 22380 9364 22389
rect 11704 22380 11756 22432
rect 56324 22380 56376 22432
rect 61752 22380 61804 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 52184 22219 52236 22228
rect 52184 22185 52193 22219
rect 52193 22185 52227 22219
rect 52227 22185 52236 22219
rect 52184 22176 52236 22185
rect 3516 22040 3568 22092
rect 7564 22083 7616 22092
rect 7564 22049 7573 22083
rect 7573 22049 7607 22083
rect 7607 22049 7616 22083
rect 7564 22040 7616 22049
rect 4620 21904 4672 21956
rect 6460 21904 6512 21956
rect 9312 22083 9364 22092
rect 9312 22049 9321 22083
rect 9321 22049 9355 22083
rect 9355 22049 9364 22083
rect 9312 22040 9364 22049
rect 9496 22083 9548 22092
rect 9496 22049 9505 22083
rect 9505 22049 9539 22083
rect 9539 22049 9548 22083
rect 9496 22040 9548 22049
rect 9772 22083 9824 22092
rect 9772 22049 9781 22083
rect 9781 22049 9815 22083
rect 9815 22049 9824 22083
rect 9772 22040 9824 22049
rect 11704 22083 11756 22092
rect 11704 22049 11713 22083
rect 11713 22049 11747 22083
rect 11747 22049 11756 22083
rect 11704 22040 11756 22049
rect 26608 22083 26660 22092
rect 4068 21836 4120 21888
rect 9772 21836 9824 21888
rect 12072 21904 12124 21956
rect 24768 21972 24820 22024
rect 26608 22049 26617 22083
rect 26617 22049 26651 22083
rect 26651 22049 26660 22083
rect 26608 22040 26660 22049
rect 35532 22040 35584 22092
rect 56324 22083 56376 22092
rect 56324 22049 56333 22083
rect 56333 22049 56367 22083
rect 56367 22049 56376 22083
rect 56324 22040 56376 22049
rect 57888 22083 57940 22092
rect 57888 22049 57897 22083
rect 57897 22049 57931 22083
rect 57931 22049 57940 22083
rect 57888 22040 57940 22049
rect 61752 22083 61804 22092
rect 61752 22049 61761 22083
rect 61761 22049 61795 22083
rect 61795 22049 61804 22083
rect 61752 22040 61804 22049
rect 26148 22015 26200 22024
rect 26148 21981 26157 22015
rect 26157 21981 26191 22015
rect 26191 21981 26200 22015
rect 26148 21972 26200 21981
rect 56324 21904 56376 21956
rect 61752 21904 61804 21956
rect 66168 21904 66220 21956
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 6460 21675 6512 21684
rect 6460 21641 6469 21675
rect 6469 21641 6503 21675
rect 6503 21641 6512 21675
rect 6460 21632 6512 21641
rect 9496 21632 9548 21684
rect 12072 21675 12124 21684
rect 12072 21641 12081 21675
rect 12081 21641 12115 21675
rect 12115 21641 12124 21675
rect 12072 21632 12124 21641
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 9680 21496 9732 21548
rect 11796 21496 11848 21548
rect 12348 21564 12400 21616
rect 26608 21632 26660 21684
rect 56324 21675 56376 21684
rect 56324 21641 56333 21675
rect 56333 21641 56367 21675
rect 56367 21641 56376 21675
rect 56324 21632 56376 21641
rect 61752 21675 61804 21684
rect 61752 21641 61761 21675
rect 61761 21641 61795 21675
rect 61795 21641 61804 21675
rect 61752 21632 61804 21641
rect 36452 21496 36504 21548
rect 56508 21496 56560 21548
rect 61660 21539 61712 21548
rect 61660 21505 61669 21539
rect 61669 21505 61703 21539
rect 61703 21505 61712 21539
rect 61660 21496 61712 21505
rect 17868 21428 17920 21480
rect 26148 21428 26200 21480
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 3976 21088 4028 21140
rect 12348 21088 12400 21140
rect 17868 20952 17920 21004
rect 8668 20884 8720 20936
rect 27160 20927 27212 20936
rect 27160 20893 27169 20927
rect 27169 20893 27203 20927
rect 27203 20893 27212 20927
rect 27160 20884 27212 20893
rect 62672 20927 62724 20936
rect 62672 20893 62681 20927
rect 62681 20893 62715 20927
rect 62715 20893 62724 20927
rect 62672 20884 62724 20893
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 8668 20451 8720 20460
rect 8668 20417 8677 20451
rect 8677 20417 8711 20451
rect 8711 20417 8720 20451
rect 8668 20408 8720 20417
rect 61660 20408 61712 20460
rect 62028 20408 62080 20460
rect 62672 20408 62724 20460
rect 64880 20451 64932 20460
rect 64880 20417 64889 20451
rect 64889 20417 64923 20451
rect 64923 20417 64932 20451
rect 64880 20408 64932 20417
rect 9036 20340 9088 20392
rect 4068 20272 4120 20324
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 9036 20043 9088 20052
rect 9036 20009 9045 20043
rect 9045 20009 9079 20043
rect 9079 20009 9088 20043
rect 9036 20000 9088 20009
rect 8392 19796 8444 19848
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 27896 19363 27948 19372
rect 27896 19329 27905 19363
rect 27905 19329 27939 19363
rect 27939 19329 27948 19363
rect 27896 19320 27948 19329
rect 34704 19320 34756 19372
rect 53380 19252 53432 19304
rect 66168 19252 66220 19304
rect 35716 19184 35768 19236
rect 27988 19159 28040 19168
rect 27988 19125 27997 19159
rect 27997 19125 28031 19159
rect 28031 19125 28040 19159
rect 27988 19116 28040 19125
rect 29000 19116 29052 19168
rect 35532 19116 35584 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 27988 18776 28040 18828
rect 29000 18819 29052 18828
rect 29000 18785 29009 18819
rect 29009 18785 29043 18819
rect 29043 18785 29052 18819
rect 29000 18776 29052 18785
rect 35532 18819 35584 18828
rect 35532 18785 35541 18819
rect 35541 18785 35575 18819
rect 35575 18785 35584 18819
rect 35532 18776 35584 18785
rect 35716 18819 35768 18828
rect 35716 18785 35725 18819
rect 35725 18785 35759 18819
rect 35759 18785 35768 18819
rect 35716 18776 35768 18785
rect 37188 18819 37240 18828
rect 37188 18785 37197 18819
rect 37197 18785 37231 18819
rect 37231 18785 37240 18819
rect 37188 18776 37240 18785
rect 24124 18708 24176 18760
rect 24768 18751 24820 18760
rect 24768 18717 24777 18751
rect 24777 18717 24811 18751
rect 24811 18717 24820 18751
rect 24768 18708 24820 18717
rect 4712 18640 4764 18692
rect 24308 18572 24360 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 24308 18343 24360 18352
rect 24308 18309 24317 18343
rect 24317 18309 24351 18343
rect 24351 18309 24360 18343
rect 24308 18300 24360 18309
rect 24124 18275 24176 18284
rect 24124 18241 24133 18275
rect 24133 18241 24167 18275
rect 24167 18241 24176 18275
rect 24124 18232 24176 18241
rect 24124 18096 24176 18148
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 52920 17824 52972 17876
rect 66168 17824 66220 17876
rect 38476 17731 38528 17740
rect 38476 17697 38485 17731
rect 38485 17697 38519 17731
rect 38519 17697 38528 17731
rect 38476 17688 38528 17697
rect 13728 17620 13780 17672
rect 33692 17620 33744 17672
rect 36820 17663 36872 17672
rect 36820 17629 36829 17663
rect 36829 17629 36863 17663
rect 36863 17629 36872 17663
rect 36820 17620 36872 17629
rect 58164 17620 58216 17672
rect 59176 17620 59228 17672
rect 59360 17484 59412 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 59360 17255 59412 17264
rect 59360 17221 59369 17255
rect 59369 17221 59403 17255
rect 59403 17221 59412 17255
rect 59360 17212 59412 17221
rect 13728 17187 13780 17196
rect 13728 17153 13737 17187
rect 13737 17153 13771 17187
rect 13771 17153 13780 17187
rect 13728 17144 13780 17153
rect 36820 17144 36872 17196
rect 59176 17187 59228 17196
rect 59176 17153 59185 17187
rect 59185 17153 59219 17187
rect 59219 17153 59228 17187
rect 59176 17144 59228 17153
rect 13912 17119 13964 17128
rect 13912 17085 13921 17119
rect 13921 17085 13955 17119
rect 13955 17085 13964 17119
rect 13912 17076 13964 17085
rect 14464 17119 14516 17128
rect 14464 17085 14473 17119
rect 14473 17085 14507 17119
rect 14507 17085 14516 17119
rect 14464 17076 14516 17085
rect 65524 17076 65576 17128
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 13912 16736 13964 16788
rect 14280 16585 14332 16594
rect 14280 16551 14289 16585
rect 14289 16551 14323 16585
rect 14323 16551 14332 16585
rect 14280 16542 14332 16551
rect 4068 16396 4120 16448
rect 4620 16396 4672 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 23112 15444 23164 15496
rect 27896 15444 27948 15496
rect 62028 15487 62080 15496
rect 62028 15453 62037 15487
rect 62037 15453 62071 15487
rect 62071 15453 62080 15487
rect 62028 15444 62080 15453
rect 62856 15487 62908 15496
rect 62856 15453 62865 15487
rect 62865 15453 62899 15487
rect 62899 15453 62908 15487
rect 62856 15444 62908 15453
rect 23756 15351 23808 15360
rect 23756 15317 23765 15351
rect 23765 15317 23799 15351
rect 23799 15317 23808 15351
rect 23756 15308 23808 15317
rect 63224 15308 63276 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 23756 15036 23808 15088
rect 63224 15079 63276 15088
rect 63224 15045 63233 15079
rect 63233 15045 63267 15079
rect 63267 15045 63276 15079
rect 63224 15036 63276 15045
rect 23112 15011 23164 15020
rect 23112 14977 23121 15011
rect 23121 14977 23155 15011
rect 23155 14977 23164 15011
rect 23112 14968 23164 14977
rect 62856 14968 62908 15020
rect 848 14832 900 14884
rect 64788 14943 64840 14952
rect 64788 14909 64797 14943
rect 64797 14909 64831 14943
rect 64831 14909 64840 14943
rect 64788 14900 64840 14909
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 14280 14356 14332 14408
rect 38844 14424 38896 14476
rect 36360 14399 36412 14408
rect 36360 14365 36369 14399
rect 36369 14365 36403 14399
rect 36403 14365 36412 14399
rect 36360 14356 36412 14365
rect 15108 14263 15160 14272
rect 15108 14229 15117 14263
rect 15117 14229 15151 14263
rect 15151 14229 15160 14263
rect 15108 14220 15160 14229
rect 35808 14263 35860 14272
rect 35808 14229 35817 14263
rect 35817 14229 35851 14263
rect 35851 14229 35860 14263
rect 35808 14220 35860 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 31944 13948 31996 14000
rect 30748 13923 30800 13932
rect 30748 13889 30757 13923
rect 30757 13889 30791 13923
rect 30791 13889 30800 13923
rect 30748 13880 30800 13889
rect 12256 13812 12308 13864
rect 32128 13812 32180 13864
rect 14924 13676 14976 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 4068 13336 4120 13388
rect 12256 13379 12308 13388
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 12256 13336 12308 13345
rect 14924 13379 14976 13388
rect 14924 13345 14933 13379
rect 14933 13345 14967 13379
rect 14967 13345 14976 13379
rect 14924 13336 14976 13345
rect 15108 13379 15160 13388
rect 15108 13345 15117 13379
rect 15117 13345 15151 13379
rect 15151 13345 15160 13379
rect 15108 13336 15160 13345
rect 15476 13379 15528 13388
rect 15476 13345 15485 13379
rect 15485 13345 15519 13379
rect 15519 13345 15528 13379
rect 15476 13336 15528 13345
rect 31944 13379 31996 13388
rect 31944 13345 31953 13379
rect 31953 13345 31987 13379
rect 31987 13345 31996 13379
rect 31944 13336 31996 13345
rect 32128 13379 32180 13388
rect 32128 13345 32137 13379
rect 32137 13345 32171 13379
rect 32171 13345 32180 13379
rect 32128 13336 32180 13345
rect 36360 13404 36412 13456
rect 35808 13379 35860 13388
rect 35808 13345 35817 13379
rect 35817 13345 35851 13379
rect 35851 13345 35860 13379
rect 35808 13336 35860 13345
rect 36084 13379 36136 13388
rect 36084 13345 36093 13379
rect 36093 13345 36127 13379
rect 36127 13345 36136 13379
rect 36084 13336 36136 13345
rect 11612 13200 11664 13252
rect 30288 13243 30340 13252
rect 30288 13209 30297 13243
rect 30297 13209 30331 13243
rect 30331 13209 30340 13243
rect 30288 13200 30340 13209
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 11612 12971 11664 12980
rect 11612 12937 11621 12971
rect 11621 12937 11655 12971
rect 11655 12937 11664 12971
rect 11612 12928 11664 12937
rect 3332 12860 3384 12912
rect 30288 12928 30340 12980
rect 11796 12792 11848 12844
rect 9036 12631 9088 12640
rect 9036 12597 9045 12631
rect 9045 12597 9079 12631
rect 9079 12597 9088 12631
rect 9036 12588 9088 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 8944 12180 8996 12232
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 40040 12180 40092 12232
rect 41512 12223 41564 12232
rect 41512 12189 41521 12223
rect 41521 12189 41555 12223
rect 41555 12189 41564 12223
rect 41512 12180 41564 12189
rect 9220 12044 9272 12096
rect 41880 12044 41932 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 9220 11815 9272 11824
rect 9220 11781 9229 11815
rect 9229 11781 9263 11815
rect 9263 11781 9272 11815
rect 9220 11772 9272 11781
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 40040 11747 40092 11756
rect 40040 11713 40049 11747
rect 40049 11713 40083 11747
rect 40083 11713 40092 11747
rect 40040 11704 40092 11713
rect 9772 11679 9824 11688
rect 9772 11645 9781 11679
rect 9781 11645 9815 11679
rect 9815 11645 9824 11679
rect 9772 11636 9824 11645
rect 40224 11679 40276 11688
rect 40224 11645 40233 11679
rect 40233 11645 40267 11679
rect 40267 11645 40276 11679
rect 40224 11636 40276 11645
rect 62120 11636 62172 11688
rect 9128 11500 9180 11552
rect 24400 11543 24452 11552
rect 24400 11509 24409 11543
rect 24409 11509 24443 11543
rect 24443 11509 24452 11543
rect 24400 11500 24452 11509
rect 41696 11500 41748 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 40224 11296 40276 11348
rect 20720 11228 20772 11280
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9128 11203 9180 11212
rect 9128 11169 9137 11203
rect 9137 11169 9171 11203
rect 9171 11169 9180 11203
rect 9128 11160 9180 11169
rect 9864 11203 9916 11212
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 9864 11160 9916 11169
rect 24400 11203 24452 11212
rect 24400 11169 24409 11203
rect 24409 11169 24443 11203
rect 24443 11169 24452 11203
rect 24400 11160 24452 11169
rect 41696 11203 41748 11212
rect 41696 11169 41705 11203
rect 41705 11169 41739 11203
rect 41739 11169 41748 11203
rect 41696 11160 41748 11169
rect 41880 11203 41932 11212
rect 41880 11169 41889 11203
rect 41889 11169 41923 11203
rect 41923 11169 41932 11203
rect 41880 11160 41932 11169
rect 27528 11135 27580 11144
rect 27528 11101 27537 11135
rect 27537 11101 27571 11135
rect 27571 11101 27580 11135
rect 27528 11092 27580 11101
rect 40132 11092 40184 11144
rect 24584 11067 24636 11076
rect 24584 11033 24593 11067
rect 24593 11033 24627 11067
rect 24627 11033 24636 11067
rect 24584 11024 24636 11033
rect 57244 11024 57296 11076
rect 3424 10956 3476 11008
rect 9772 10956 9824 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 24584 10752 24636 10804
rect 9680 10616 9732 10668
rect 24860 10659 24912 10668
rect 24860 10625 24869 10659
rect 24869 10625 24903 10659
rect 24903 10625 24912 10659
rect 24860 10616 24912 10625
rect 27528 10659 27580 10668
rect 27528 10625 27537 10659
rect 27537 10625 27571 10659
rect 27571 10625 27580 10659
rect 27528 10616 27580 10625
rect 38200 10659 38252 10668
rect 38200 10625 38209 10659
rect 38209 10625 38243 10659
rect 38243 10625 38252 10659
rect 38200 10616 38252 10625
rect 40132 10616 40184 10668
rect 62120 10616 62172 10668
rect 66168 10616 66220 10668
rect 27896 10548 27948 10600
rect 29368 10591 29420 10600
rect 29368 10557 29377 10591
rect 29377 10557 29411 10591
rect 29411 10557 29420 10591
rect 29368 10548 29420 10557
rect 9772 10412 9824 10464
rect 9956 10412 10008 10464
rect 38292 10455 38344 10464
rect 38292 10421 38301 10455
rect 38301 10421 38335 10455
rect 38335 10421 38344 10455
rect 38292 10412 38344 10421
rect 38844 10455 38896 10464
rect 38844 10421 38853 10455
rect 38853 10421 38887 10455
rect 38887 10421 38896 10455
rect 38844 10412 38896 10421
rect 44088 10455 44140 10464
rect 44088 10421 44097 10455
rect 44097 10421 44131 10455
rect 44131 10421 44140 10455
rect 44088 10412 44140 10421
rect 45008 10412 45060 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 27896 10251 27948 10260
rect 27896 10217 27905 10251
rect 27905 10217 27939 10251
rect 27939 10217 27948 10251
rect 27896 10208 27948 10217
rect 44088 10140 44140 10192
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 9956 10115 10008 10124
rect 9956 10081 9965 10115
rect 9965 10081 9999 10115
rect 9999 10081 10008 10115
rect 9956 10072 10008 10081
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 45008 10115 45060 10124
rect 45008 10081 45017 10115
rect 45017 10081 45051 10115
rect 45051 10081 45060 10115
rect 45008 10072 45060 10081
rect 24860 10004 24912 10056
rect 38200 10004 38252 10056
rect 62764 9936 62816 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 3424 9596 3476 9648
rect 9864 9596 9916 9648
rect 38292 9639 38344 9648
rect 38292 9605 38301 9639
rect 38301 9605 38335 9639
rect 38335 9605 38344 9639
rect 38292 9596 38344 9605
rect 38660 9503 38712 9512
rect 38660 9469 38669 9503
rect 38669 9469 38703 9503
rect 38703 9469 38712 9503
rect 38660 9460 38712 9469
rect 38844 9392 38896 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 3424 8236 3476 8288
rect 20720 8236 20772 8288
rect 47768 8236 47820 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 47768 7939 47820 7948
rect 47768 7905 47777 7939
rect 47777 7905 47811 7939
rect 47811 7905 47820 7939
rect 47768 7896 47820 7905
rect 47124 7871 47176 7880
rect 47124 7837 47133 7871
rect 47133 7837 47167 7871
rect 47167 7837 47176 7871
rect 47124 7828 47176 7837
rect 66168 7760 66220 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 43260 6808 43312 6860
rect 47124 6808 47176 6860
rect 11152 6740 11204 6792
rect 10784 6672 10836 6724
rect 10968 6672 11020 6724
rect 11520 6740 11572 6792
rect 11704 6604 11756 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 11704 6375 11756 6384
rect 11704 6341 11713 6375
rect 11713 6341 11747 6375
rect 11747 6341 11756 6375
rect 11704 6332 11756 6341
rect 10784 6307 10836 6316
rect 10784 6273 10793 6307
rect 10793 6273 10827 6307
rect 10827 6273 10836 6307
rect 10784 6264 10836 6273
rect 11520 6307 11572 6316
rect 11520 6273 11529 6307
rect 11529 6273 11563 6307
rect 11563 6273 11572 6307
rect 11520 6264 11572 6273
rect 43260 6264 43312 6316
rect 12440 6239 12492 6248
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 12440 6196 12492 6205
rect 11336 6060 11388 6112
rect 43628 6060 43680 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 9036 5788 9088 5840
rect 11152 5763 11204 5772
rect 11152 5729 11161 5763
rect 11161 5729 11195 5763
rect 11195 5729 11204 5763
rect 11152 5720 11204 5729
rect 11336 5763 11388 5772
rect 11336 5729 11345 5763
rect 11345 5729 11379 5763
rect 11379 5729 11388 5763
rect 11336 5720 11388 5729
rect 43444 5652 43496 5704
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 3424 5312 3476 5364
rect 12440 5312 12492 5364
rect 3148 5244 3200 5296
rect 10324 5244 10376 5296
rect 43628 5287 43680 5296
rect 43628 5253 43637 5287
rect 43637 5253 43671 5287
rect 43671 5253 43680 5287
rect 43628 5244 43680 5253
rect 43444 5219 43496 5228
rect 43444 5185 43453 5219
rect 43453 5185 43487 5219
rect 43487 5185 43496 5219
rect 43444 5176 43496 5185
rect 60648 5108 60700 5160
rect 13544 4972 13596 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 29000 4700 29052 4752
rect 13544 4675 13596 4684
rect 13544 4641 13553 4675
rect 13553 4641 13587 4675
rect 13587 4641 13596 4675
rect 13544 4632 13596 4641
rect 29552 4564 29604 4616
rect 11612 4496 11664 4548
rect 13360 4539 13412 4548
rect 13360 4505 13369 4539
rect 13369 4505 13403 4539
rect 13403 4505 13412 4539
rect 13360 4496 13412 4505
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 13360 4224 13412 4276
rect 11796 4088 11848 4140
rect 28816 4088 28868 4140
rect 29000 4131 29052 4140
rect 29000 4097 29009 4131
rect 29009 4097 29043 4131
rect 29043 4097 29052 4131
rect 29000 4088 29052 4097
rect 62764 4088 62816 4140
rect 66168 4088 66220 4140
rect 29644 4063 29696 4072
rect 29644 4029 29653 4063
rect 29653 4029 29687 4063
rect 29687 4029 29696 4063
rect 29644 4020 29696 4029
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 54576 3612 54628 3664
rect 67640 3612 67692 3664
rect 24492 3544 24544 3596
rect 29368 3544 29420 3596
rect 29552 3587 29604 3596
rect 29552 3553 29561 3587
rect 29561 3553 29595 3587
rect 29595 3553 29604 3587
rect 29552 3544 29604 3553
rect 56048 3544 56100 3596
rect 57336 3544 57388 3596
rect 57612 3544 57664 3596
rect 58624 3544 58676 3596
rect 6460 3476 6512 3528
rect 14464 3476 14516 3528
rect 18052 3476 18104 3528
rect 24124 3476 24176 3528
rect 28816 3519 28868 3528
rect 28816 3485 28825 3519
rect 28825 3485 28859 3519
rect 28859 3485 28868 3519
rect 28816 3476 28868 3485
rect 37188 3476 37240 3528
rect 68928 3476 68980 3528
rect 10324 3408 10376 3460
rect 24676 3408 24728 3460
rect 65064 3408 65116 3460
rect 57888 3340 57940 3392
rect 59912 3340 59964 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 60648 2796 60700 2848
rect 63776 2796 63828 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
<< metal2 >>
rect 634 71200 746 72000
rect 1922 71200 2034 72000
rect 3210 71200 3322 72000
rect 4498 71200 4610 72000
rect 5786 71200 5898 72000
rect 7074 71200 7186 72000
rect 8362 71200 8474 72000
rect 9650 71200 9762 72000
rect 10938 71200 11050 72000
rect 12226 71200 12338 72000
rect 13514 71200 13626 72000
rect 14802 71200 14914 72000
rect 16090 71200 16202 72000
rect 17378 71200 17490 72000
rect 18666 71200 18778 72000
rect 19954 71200 20066 72000
rect 21242 71200 21354 72000
rect 22530 71200 22642 72000
rect 24462 71200 24574 72000
rect 25750 71200 25862 72000
rect 27038 71200 27150 72000
rect 28326 71200 28438 72000
rect 29614 71200 29726 72000
rect 30902 71200 31014 72000
rect 32190 71346 32302 72000
rect 31772 71318 32302 71346
rect 1964 68338 1992 71200
rect 1952 68332 2004 68338
rect 1952 68274 2004 68280
rect 1400 66156 1452 66162
rect 1400 66098 1452 66104
rect 1412 66065 1440 66098
rect 1584 66088 1636 66094
rect 1398 66056 1454 66065
rect 1584 66030 1636 66036
rect 1398 65991 1454 66000
rect 1596 36854 1624 66030
rect 3252 64874 3280 71200
rect 4214 69116 4522 69136
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69040 4522 69060
rect 3606 68776 3662 68785
rect 3606 68711 3662 68720
rect 3514 67416 3570 67425
rect 3514 67351 3570 67360
rect 2792 64846 3280 64874
rect 2792 56302 2820 64846
rect 3330 64696 3386 64705
rect 3330 64631 3386 64640
rect 3344 60602 3372 64631
rect 3422 61976 3478 61985
rect 3422 61911 3478 61920
rect 3436 60790 3464 61911
rect 3424 60784 3476 60790
rect 3424 60726 3476 60732
rect 3344 60574 3464 60602
rect 3330 59256 3386 59265
rect 3330 59191 3386 59200
rect 2780 56296 2832 56302
rect 2780 56238 2832 56244
rect 3344 55282 3372 59191
rect 3332 55276 3384 55282
rect 3332 55218 3384 55224
rect 1584 36848 1636 36854
rect 1584 36790 1636 36796
rect 3436 34218 3464 60574
rect 3528 35894 3556 67351
rect 3620 39370 3648 68711
rect 4214 68028 4522 68048
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67952 4522 67972
rect 4214 66940 4522 66960
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66864 4522 66884
rect 4214 65852 4522 65872
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65776 4522 65796
rect 5828 64874 5856 71200
rect 7116 64874 7144 71200
rect 14844 64874 14872 71200
rect 15844 68332 15896 68338
rect 15844 68274 15896 68280
rect 5552 64846 5856 64874
rect 6932 64846 7144 64874
rect 13832 64846 14872 64874
rect 4214 64764 4522 64784
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64688 4522 64708
rect 4214 63676 4522 63696
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63600 4522 63620
rect 4214 62588 4522 62608
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62512 4522 62532
rect 5552 62218 5580 64846
rect 5540 62212 5592 62218
rect 5540 62154 5592 62160
rect 4214 61500 4522 61520
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61424 4522 61444
rect 4214 60412 4522 60432
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60336 4522 60356
rect 4214 59324 4522 59344
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59248 4522 59268
rect 4214 58236 4522 58256
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58160 4522 58180
rect 3698 57896 3754 57905
rect 3698 57831 3754 57840
rect 3712 48074 3740 57831
rect 4214 57148 4522 57168
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57072 4522 57092
rect 4214 56060 4522 56080
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55984 4522 56004
rect 4214 54972 4522 54992
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54896 4522 54916
rect 4214 53884 4522 53904
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53808 4522 53828
rect 4214 52796 4522 52816
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52720 4522 52740
rect 4214 51708 4522 51728
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51632 4522 51652
rect 4214 50620 4522 50640
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50544 4522 50564
rect 6932 50386 6960 64846
rect 6920 50380 6972 50386
rect 6920 50322 6972 50328
rect 4214 49532 4522 49552
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49456 4522 49476
rect 4214 48444 4522 48464
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48368 4522 48388
rect 3700 48068 3752 48074
rect 3700 48010 3752 48016
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 3698 46336 3754 46345
rect 3698 46271 3754 46280
rect 3712 42770 3740 46271
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 3700 42764 3752 42770
rect 3700 42706 3752 42712
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 9772 39840 9824 39846
rect 9772 39782 9824 39788
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 9784 39506 9812 39782
rect 9772 39500 9824 39506
rect 9772 39442 9824 39448
rect 3608 39364 3660 39370
rect 3608 39306 3660 39312
rect 10416 39364 10468 39370
rect 10416 39306 10468 39312
rect 10428 39098 10456 39306
rect 10416 39092 10468 39098
rect 10416 39034 10468 39040
rect 10508 38956 10560 38962
rect 10508 38898 10560 38904
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 6368 36168 6420 36174
rect 6368 36110 6420 36116
rect 3528 35866 3648 35894
rect 3436 34190 3556 34218
rect 3422 34096 3478 34105
rect 3422 34031 3478 34040
rect 3436 33930 3464 34031
rect 3424 33924 3476 33930
rect 3424 33866 3476 33872
rect 2962 31376 3018 31385
rect 2962 31311 3018 31320
rect 2976 30870 3004 31311
rect 2964 30864 3016 30870
rect 2964 30806 3016 30812
rect 3424 28960 3476 28966
rect 3424 28902 3476 28908
rect 3436 28665 3464 28902
rect 3422 28656 3478 28665
rect 3422 28591 3478 28600
rect 3146 25936 3202 25945
rect 3146 25871 3202 25880
rect 3160 25226 3188 25871
rect 3148 25220 3200 25226
rect 3148 25162 3200 25168
rect 3424 24676 3476 24682
rect 3424 24618 3476 24624
rect 3436 24585 3464 24618
rect 3422 24576 3478 24585
rect 3422 24511 3478 24520
rect 3528 22098 3556 34190
rect 3620 30122 3648 35866
rect 6380 35698 6408 36110
rect 6368 35692 6420 35698
rect 6368 35634 6420 35640
rect 6552 35624 6604 35630
rect 6552 35566 6604 35572
rect 4068 35556 4120 35562
rect 4068 35498 4120 35504
rect 4080 35465 4108 35498
rect 4066 35456 4122 35465
rect 4066 35391 4122 35400
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 6564 35290 6592 35566
rect 6552 35284 6604 35290
rect 6552 35226 6604 35232
rect 6552 35080 6604 35086
rect 6552 35022 6604 35028
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 5460 30802 5488 31758
rect 6564 31346 6592 35022
rect 10520 34542 10548 38898
rect 13832 36650 13860 64846
rect 15856 63510 15884 68274
rect 17420 64874 17448 71200
rect 18708 64874 18736 71200
rect 19574 69660 19882 69680
rect 19574 69658 19580 69660
rect 19636 69658 19660 69660
rect 19716 69658 19740 69660
rect 19796 69658 19820 69660
rect 19876 69658 19882 69660
rect 19636 69606 19638 69658
rect 19818 69606 19820 69658
rect 19574 69604 19580 69606
rect 19636 69604 19660 69606
rect 19716 69604 19740 69606
rect 19796 69604 19820 69606
rect 19876 69604 19882 69606
rect 19574 69584 19882 69604
rect 19574 68572 19882 68592
rect 19574 68570 19580 68572
rect 19636 68570 19660 68572
rect 19716 68570 19740 68572
rect 19796 68570 19820 68572
rect 19876 68570 19882 68572
rect 19636 68518 19638 68570
rect 19818 68518 19820 68570
rect 19574 68516 19580 68518
rect 19636 68516 19660 68518
rect 19716 68516 19740 68518
rect 19796 68516 19820 68518
rect 19876 68516 19882 68518
rect 19574 68496 19882 68516
rect 19996 67794 20024 71200
rect 21284 68338 21312 71200
rect 21272 68332 21324 68338
rect 21272 68274 21324 68280
rect 19984 67788 20036 67794
rect 19984 67730 20036 67736
rect 21272 67788 21324 67794
rect 21272 67730 21324 67736
rect 19574 67484 19882 67504
rect 19574 67482 19580 67484
rect 19636 67482 19660 67484
rect 19716 67482 19740 67484
rect 19796 67482 19820 67484
rect 19876 67482 19882 67484
rect 19636 67430 19638 67482
rect 19818 67430 19820 67482
rect 19574 67428 19580 67430
rect 19636 67428 19660 67430
rect 19716 67428 19740 67430
rect 19796 67428 19820 67430
rect 19876 67428 19882 67430
rect 19574 67408 19882 67428
rect 19574 66396 19882 66416
rect 19574 66394 19580 66396
rect 19636 66394 19660 66396
rect 19716 66394 19740 66396
rect 19796 66394 19820 66396
rect 19876 66394 19882 66396
rect 19636 66342 19638 66394
rect 19818 66342 19820 66394
rect 19574 66340 19580 66342
rect 19636 66340 19660 66342
rect 19716 66340 19740 66342
rect 19796 66340 19820 66342
rect 19876 66340 19882 66342
rect 19574 66320 19882 66340
rect 19574 65308 19882 65328
rect 19574 65306 19580 65308
rect 19636 65306 19660 65308
rect 19716 65306 19740 65308
rect 19796 65306 19820 65308
rect 19876 65306 19882 65308
rect 19636 65254 19638 65306
rect 19818 65254 19820 65306
rect 19574 65252 19580 65254
rect 19636 65252 19660 65254
rect 19716 65252 19740 65254
rect 19796 65252 19820 65254
rect 19876 65252 19882 65254
rect 19574 65232 19882 65252
rect 16592 64846 17448 64874
rect 17972 64846 18736 64874
rect 15844 63504 15896 63510
rect 15844 63446 15896 63452
rect 16592 42566 16620 64846
rect 16764 43104 16816 43110
rect 16764 43046 16816 43052
rect 16776 42702 16804 43046
rect 16764 42696 16816 42702
rect 16764 42638 16816 42644
rect 16948 42628 17000 42634
rect 16948 42570 17000 42576
rect 16580 42560 16632 42566
rect 16580 42502 16632 42508
rect 16960 42362 16988 42570
rect 16948 42356 17000 42362
rect 16948 42298 17000 42304
rect 14464 42220 14516 42226
rect 14464 42162 14516 42168
rect 14188 36712 14240 36718
rect 14188 36654 14240 36660
rect 13820 36644 13872 36650
rect 13820 36586 13872 36592
rect 14200 36378 14228 36654
rect 14188 36372 14240 36378
rect 14188 36314 14240 36320
rect 14280 36168 14332 36174
rect 14280 36110 14332 36116
rect 14292 35630 14320 36110
rect 14280 35624 14332 35630
rect 14280 35566 14332 35572
rect 14292 35086 14320 35566
rect 14280 35080 14332 35086
rect 14280 35022 14332 35028
rect 10508 34536 10560 34542
rect 10508 34478 10560 34484
rect 10968 34536 11020 34542
rect 10968 34478 11020 34484
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 5632 31136 5684 31142
rect 5632 31078 5684 31084
rect 5644 30802 5672 31078
rect 5448 30796 5500 30802
rect 5448 30738 5500 30744
rect 5632 30796 5684 30802
rect 5632 30738 5684 30744
rect 3608 30116 3660 30122
rect 3608 30058 3660 30064
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3516 22092 3568 22098
rect 3516 22034 3568 22040
rect 848 14884 900 14890
rect 848 14826 900 14832
rect -10 0 102 800
rect 860 762 888 14826
rect 3332 12912 3384 12918
rect 3332 12854 3384 12860
rect 3344 6914 3372 12854
rect 3620 12434 3648 24550
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4620 21956 4672 21962
rect 4620 21898 4672 21904
rect 6460 21956 6512 21962
rect 6460 21898 6512 21904
rect 4068 21888 4120 21894
rect 4066 21856 4068 21865
rect 4120 21856 4122 21865
rect 4066 21791 4122 21800
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 3988 15065 4016 21082
rect 4066 20496 4122 20505
rect 4066 20431 4122 20440
rect 4080 20330 4108 20431
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4632 16454 4660 21898
rect 6472 21690 6500 21898
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6564 21554 6592 31282
rect 7748 30728 7800 30734
rect 7748 30670 7800 30676
rect 7760 30258 7788 30670
rect 7748 30252 7800 30258
rect 7748 30194 7800 30200
rect 8300 30184 8352 30190
rect 8300 30126 8352 30132
rect 8312 29850 8340 30126
rect 8300 29844 8352 29850
rect 8300 29786 8352 29792
rect 8392 29640 8444 29646
rect 8392 29582 8444 29588
rect 8404 28490 8432 29582
rect 8392 28484 8444 28490
rect 8392 28426 8444 28432
rect 9128 28484 9180 28490
rect 9128 28426 9180 28432
rect 6920 26852 6972 26858
rect 6920 26794 6972 26800
rect 6932 22094 6960 26794
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 7576 22098 7604 22374
rect 6932 22066 7328 22094
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4068 16448 4120 16454
rect 4066 16416 4068 16425
rect 4620 16448 4672 16454
rect 4120 16416 4122 16425
rect 4620 16390 4672 16396
rect 4066 16351 4122 16360
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 3974 15056 4030 15065
rect 3974 14991 4030 15000
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4066 13696 4122 13705
rect 4066 13631 4122 13640
rect 4080 13394 4108 13631
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 3528 12406 3648 12434
rect 3424 11008 3476 11014
rect 3422 10976 3424 10985
rect 3476 10976 3478 10985
rect 3422 10911 3478 10920
rect 3424 9648 3476 9654
rect 3422 9616 3424 9625
rect 3476 9616 3478 9625
rect 3422 9551 3478 9560
rect 3424 8288 3476 8294
rect 3422 8256 3424 8265
rect 3476 8256 3478 8265
rect 3422 8191 3478 8200
rect 3344 6905 3464 6914
rect 3344 6896 3478 6905
rect 3344 6886 3422 6896
rect 3422 6831 3478 6840
rect 3422 5536 3478 5545
rect 3422 5471 3478 5480
rect 3436 5370 3464 5471
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 3160 4185 3188 5238
rect 3146 4176 3202 4185
rect 3146 4111 3202 4120
rect 3528 2825 3556 12406
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3514 2816 3570 2825
rect 3514 2751 3570 2760
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 1136 870 1348 898
rect 1136 762 1164 870
rect 1320 800 1348 870
rect 860 734 1164 762
rect 1278 0 1390 800
rect 2566 0 2678 800
rect 3854 0 3966 800
rect 4724 762 4752 18634
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5000 870 5212 898
rect 5000 762 5028 870
rect 5184 800 5212 870
rect 6472 800 6500 3470
rect 4724 734 5028 762
rect 5142 0 5254 800
rect 6430 0 6542 800
rect 7300 762 7328 22066
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8680 20466 8708 20878
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9048 20058 9076 20334
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9140 19854 9168 28426
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9324 22098 9352 22374
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9496 22092 9548 22098
rect 9496 22034 9548 22040
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9508 21690 9536 22034
rect 9784 21894 9812 22034
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8404 11762 8432 19790
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8956 11218 8984 12174
rect 9048 11762 9076 12582
rect 9692 12238 9720 21490
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9232 11830 9260 12038
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9140 11218 9168 11494
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9692 10674 9720 12174
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9784 11014 9812 11630
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10130 9812 10406
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9876 9654 9904 11154
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 10130 9996 10406
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 7576 870 7788 898
rect 7576 762 7604 870
rect 7760 800 7788 870
rect 9048 800 9076 5782
rect 10336 5302 10364 10066
rect 10980 6730 11008 34478
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12360 24818 12388 25230
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12992 24744 13044 24750
rect 12992 24686 13044 24692
rect 13004 24410 13032 24686
rect 12992 24404 13044 24410
rect 12992 24346 13044 24352
rect 14476 24206 14504 42162
rect 17972 29238 18000 64846
rect 19432 64456 19484 64462
rect 19432 64398 19484 64404
rect 19444 63986 19472 64398
rect 19574 64220 19882 64240
rect 19574 64218 19580 64220
rect 19636 64218 19660 64220
rect 19716 64218 19740 64220
rect 19796 64218 19820 64220
rect 19876 64218 19882 64220
rect 19636 64166 19638 64218
rect 19818 64166 19820 64218
rect 19574 64164 19580 64166
rect 19636 64164 19660 64166
rect 19716 64164 19740 64166
rect 19796 64164 19820 64166
rect 19876 64164 19882 64166
rect 19574 64144 19882 64164
rect 21284 64054 21312 67730
rect 21272 64048 21324 64054
rect 21272 63990 21324 63996
rect 19432 63980 19484 63986
rect 19432 63922 19484 63928
rect 20168 63912 20220 63918
rect 20168 63854 20220 63860
rect 19340 63776 19392 63782
rect 19340 63718 19392 63724
rect 19352 63442 19380 63718
rect 19340 63436 19392 63442
rect 19340 63378 19392 63384
rect 19432 63232 19484 63238
rect 19432 63174 19484 63180
rect 19444 63034 19472 63174
rect 19574 63132 19882 63152
rect 19574 63130 19580 63132
rect 19636 63130 19660 63132
rect 19716 63130 19740 63132
rect 19796 63130 19820 63132
rect 19876 63130 19882 63132
rect 19636 63078 19638 63130
rect 19818 63078 19820 63130
rect 19574 63076 19580 63078
rect 19636 63076 19660 63078
rect 19716 63076 19740 63078
rect 19796 63076 19820 63078
rect 19876 63076 19882 63078
rect 19574 63056 19882 63076
rect 20180 63034 20208 63854
rect 19432 63028 19484 63034
rect 19432 62970 19484 62976
rect 20168 63028 20220 63034
rect 20168 62970 20220 62976
rect 19574 62044 19882 62064
rect 19574 62042 19580 62044
rect 19636 62042 19660 62044
rect 19716 62042 19740 62044
rect 19796 62042 19820 62044
rect 19876 62042 19882 62044
rect 19636 61990 19638 62042
rect 19818 61990 19820 62042
rect 19574 61988 19580 61990
rect 19636 61988 19660 61990
rect 19716 61988 19740 61990
rect 19796 61988 19820 61990
rect 19876 61988 19882 61990
rect 19574 61968 19882 61988
rect 19574 60956 19882 60976
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60880 19882 60900
rect 24860 60784 24912 60790
rect 24860 60726 24912 60732
rect 19574 59868 19882 59888
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59792 19882 59812
rect 24872 59498 24900 60726
rect 26976 60104 27028 60110
rect 26976 60046 27028 60052
rect 26988 59634 27016 60046
rect 26240 59628 26292 59634
rect 26240 59570 26292 59576
rect 26976 59628 27028 59634
rect 26976 59570 27028 59576
rect 24860 59492 24912 59498
rect 24860 59434 24912 59440
rect 19574 58780 19882 58800
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58704 19882 58724
rect 19574 57692 19882 57712
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57616 19882 57636
rect 19574 56604 19882 56624
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56528 19882 56548
rect 19574 55516 19882 55536
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55440 19882 55460
rect 19574 54428 19882 54448
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54352 19882 54372
rect 19574 53340 19882 53360
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53264 19882 53284
rect 19574 52252 19882 52272
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52176 19882 52196
rect 19574 51164 19882 51184
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51088 19882 51108
rect 24400 50720 24452 50726
rect 24400 50662 24452 50668
rect 24412 50318 24440 50662
rect 24400 50312 24452 50318
rect 24400 50254 24452 50260
rect 24860 50244 24912 50250
rect 24860 50186 24912 50192
rect 19574 50076 19882 50096
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50000 19882 50020
rect 24872 49978 24900 50186
rect 24860 49972 24912 49978
rect 24860 49914 24912 49920
rect 19574 48988 19882 49008
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48912 19882 48932
rect 22652 48544 22704 48550
rect 22652 48486 22704 48492
rect 22664 48210 22692 48486
rect 22652 48204 22704 48210
rect 22652 48146 22704 48152
rect 21916 48068 21968 48074
rect 21916 48010 21968 48016
rect 19574 47900 19882 47920
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47824 19882 47844
rect 21928 47802 21956 48010
rect 21916 47796 21968 47802
rect 21916 47738 21968 47744
rect 22008 47660 22060 47666
rect 22008 47602 22060 47608
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 22020 34474 22048 47602
rect 25320 36304 25372 36310
rect 25320 36246 25372 36252
rect 25332 34474 25360 36246
rect 26252 36038 26280 59570
rect 31772 51882 31800 71318
rect 32190 71200 32302 71318
rect 33478 71200 33590 72000
rect 34766 71200 34878 72000
rect 36054 71200 36166 72000
rect 37342 71200 37454 72000
rect 38630 71200 38742 72000
rect 39918 71200 40030 72000
rect 41206 71346 41318 72000
rect 42494 71346 42606 72000
rect 40144 71318 41318 71346
rect 34808 68490 34836 71200
rect 34934 69116 35242 69136
rect 34934 69114 34940 69116
rect 34996 69114 35020 69116
rect 35076 69114 35100 69116
rect 35156 69114 35180 69116
rect 35236 69114 35242 69116
rect 34996 69062 34998 69114
rect 35178 69062 35180 69114
rect 34934 69060 34940 69062
rect 34996 69060 35020 69062
rect 35076 69060 35100 69062
rect 35156 69060 35180 69062
rect 35236 69060 35242 69062
rect 34934 69040 35242 69060
rect 34808 68462 35848 68490
rect 35348 68332 35400 68338
rect 35348 68274 35400 68280
rect 34934 68028 35242 68048
rect 34934 68026 34940 68028
rect 34996 68026 35020 68028
rect 35076 68026 35100 68028
rect 35156 68026 35180 68028
rect 35236 68026 35242 68028
rect 34996 67974 34998 68026
rect 35178 67974 35180 68026
rect 34934 67972 34940 67974
rect 34996 67972 35020 67974
rect 35076 67972 35100 67974
rect 35156 67972 35180 67974
rect 35236 67972 35242 67974
rect 34934 67952 35242 67972
rect 34934 66940 35242 66960
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66864 35242 66884
rect 34934 65852 35242 65872
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65776 35242 65796
rect 34934 64764 35242 64784
rect 34934 64762 34940 64764
rect 34996 64762 35020 64764
rect 35076 64762 35100 64764
rect 35156 64762 35180 64764
rect 35236 64762 35242 64764
rect 34996 64710 34998 64762
rect 35178 64710 35180 64762
rect 34934 64708 34940 64710
rect 34996 64708 35020 64710
rect 35076 64708 35100 64710
rect 35156 64708 35180 64710
rect 35236 64708 35242 64710
rect 34934 64688 35242 64708
rect 34934 63676 35242 63696
rect 34934 63674 34940 63676
rect 34996 63674 35020 63676
rect 35076 63674 35100 63676
rect 35156 63674 35180 63676
rect 35236 63674 35242 63676
rect 34996 63622 34998 63674
rect 35178 63622 35180 63674
rect 34934 63620 34940 63622
rect 34996 63620 35020 63622
rect 35076 63620 35100 63622
rect 35156 63620 35180 63622
rect 35236 63620 35242 63622
rect 34934 63600 35242 63620
rect 34934 62588 35242 62608
rect 34934 62586 34940 62588
rect 34996 62586 35020 62588
rect 35076 62586 35100 62588
rect 35156 62586 35180 62588
rect 35236 62586 35242 62588
rect 34996 62534 34998 62586
rect 35178 62534 35180 62586
rect 34934 62532 34940 62534
rect 34996 62532 35020 62534
rect 35076 62532 35100 62534
rect 35156 62532 35180 62534
rect 35236 62532 35242 62534
rect 34934 62512 35242 62532
rect 32772 62280 32824 62286
rect 32772 62222 32824 62228
rect 32588 62212 32640 62218
rect 32588 62154 32640 62160
rect 32600 61946 32628 62154
rect 32588 61940 32640 61946
rect 32588 61882 32640 61888
rect 32784 61742 32812 62222
rect 32772 61736 32824 61742
rect 32772 61678 32824 61684
rect 34934 61500 35242 61520
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61424 35242 61444
rect 34934 60412 35242 60432
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60336 35242 60356
rect 34934 59324 35242 59344
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59248 35242 59268
rect 34934 58236 35242 58256
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58160 35242 58180
rect 35360 57934 35388 68274
rect 35624 61804 35676 61810
rect 35624 61746 35676 61752
rect 35532 60104 35584 60110
rect 35532 60046 35584 60052
rect 35544 59090 35572 60046
rect 35532 59084 35584 59090
rect 35532 59026 35584 59032
rect 35636 58562 35664 61746
rect 35716 58948 35768 58954
rect 35716 58890 35768 58896
rect 35728 58682 35756 58890
rect 35716 58676 35768 58682
rect 35716 58618 35768 58624
rect 35440 58540 35492 58546
rect 35636 58534 35756 58562
rect 35440 58482 35492 58488
rect 34704 57928 34756 57934
rect 34704 57870 34756 57876
rect 35348 57928 35400 57934
rect 35348 57870 35400 57876
rect 34716 57526 34744 57870
rect 34704 57520 34756 57526
rect 34704 57462 34756 57468
rect 34428 57384 34480 57390
rect 34428 57326 34480 57332
rect 34440 57050 34468 57326
rect 34934 57148 35242 57168
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57072 35242 57092
rect 34428 57044 34480 57050
rect 34428 56986 34480 56992
rect 35452 56846 35480 58482
rect 35440 56840 35492 56846
rect 35440 56782 35492 56788
rect 32956 56296 33008 56302
rect 32956 56238 33008 56244
rect 33140 56296 33192 56302
rect 33140 56238 33192 56244
rect 32968 55962 32996 56238
rect 32956 55956 33008 55962
rect 32956 55898 33008 55904
rect 33152 54874 33180 56238
rect 34934 56060 35242 56080
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55984 35242 56004
rect 35452 55758 35480 56782
rect 35348 55752 35400 55758
rect 35348 55694 35400 55700
rect 35440 55752 35492 55758
rect 35440 55694 35492 55700
rect 35360 55282 35388 55694
rect 35348 55276 35400 55282
rect 35348 55218 35400 55224
rect 34796 55208 34848 55214
rect 34796 55150 34848 55156
rect 34808 54874 34836 55150
rect 34934 54972 35242 54992
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54896 35242 54916
rect 33140 54868 33192 54874
rect 33140 54810 33192 54816
rect 34796 54868 34848 54874
rect 34796 54810 34848 54816
rect 34934 53884 35242 53904
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53808 35242 53828
rect 34934 52796 35242 52816
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52720 35242 52740
rect 32312 51944 32364 51950
rect 32312 51886 32364 51892
rect 31760 51876 31812 51882
rect 31760 51818 31812 51824
rect 32324 51610 32352 51886
rect 34934 51708 35242 51728
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51632 35242 51652
rect 32312 51604 32364 51610
rect 32312 51546 32364 51552
rect 34934 50620 35242 50640
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50544 35242 50564
rect 35348 49836 35400 49842
rect 35348 49778 35400 49784
rect 34934 49532 35242 49552
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49456 35242 49476
rect 34934 48444 35242 48464
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48368 35242 48388
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34704 43104 34756 43110
rect 34704 43046 34756 43052
rect 34716 42702 34744 43046
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34704 42696 34756 42702
rect 34704 42638 34756 42644
rect 34612 42628 34664 42634
rect 34612 42570 34664 42576
rect 34624 42362 34652 42570
rect 34612 42356 34664 42362
rect 34612 42298 34664 42304
rect 32864 42220 32916 42226
rect 32864 42162 32916 42168
rect 32876 38350 32904 42162
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 32956 39432 33008 39438
rect 32956 39374 33008 39380
rect 32968 38962 32996 39374
rect 32956 38956 33008 38962
rect 32956 38898 33008 38904
rect 33140 38888 33192 38894
rect 33140 38830 33192 38836
rect 33152 38554 33180 38830
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 33140 38548 33192 38554
rect 33140 38490 33192 38496
rect 32864 38344 32916 38350
rect 32864 38286 32916 38292
rect 32404 37188 32456 37194
rect 32404 37130 32456 37136
rect 32416 36854 32444 37130
rect 32496 37120 32548 37126
rect 32496 37062 32548 37068
rect 32508 36854 32536 37062
rect 32404 36848 32456 36854
rect 32404 36790 32456 36796
rect 32496 36848 32548 36854
rect 32496 36790 32548 36796
rect 32508 36174 32536 36790
rect 32496 36168 32548 36174
rect 32496 36110 32548 36116
rect 26240 36032 26292 36038
rect 26240 35974 26292 35980
rect 32508 35698 32536 36110
rect 32772 36100 32824 36106
rect 32772 36042 32824 36048
rect 32496 35692 32548 35698
rect 32496 35634 32548 35640
rect 22008 34468 22060 34474
rect 22008 34410 22060 34416
rect 25320 34468 25372 34474
rect 25320 34410 25372 34416
rect 24860 34400 24912 34406
rect 24860 34342 24912 34348
rect 24872 34066 24900 34342
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 25228 33924 25280 33930
rect 25228 33866 25280 33872
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 25240 33658 25268 33866
rect 25228 33652 25280 33658
rect 25228 33594 25280 33600
rect 25332 33522 25360 34410
rect 25320 33516 25372 33522
rect 25320 33458 25372 33464
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 27988 30728 28040 30734
rect 27988 30670 28040 30676
rect 19444 30258 19472 30670
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 28000 30258 28028 30670
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 27804 30252 27856 30258
rect 27804 30194 27856 30200
rect 27988 30252 28040 30258
rect 27988 30194 28040 30200
rect 19984 30184 20036 30190
rect 19984 30126 20036 30132
rect 19340 30116 19392 30122
rect 19340 30058 19392 30064
rect 17960 29232 18012 29238
rect 17960 29174 18012 29180
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 11716 22098 11744 22374
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 12084 21690 12112 21898
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11624 12986 11652 13194
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11808 12850 11836 21490
rect 12360 21146 12388 21558
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13740 17202 13768 17614
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13924 16794 13952 17070
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 14292 16600 14320 24142
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17880 21010 17908 21422
rect 17868 21004 17920 21010
rect 17868 20946 17920 20952
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14280 16594 14332 16600
rect 14280 16536 14332 16542
rect 14292 14414 14320 16536
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12268 13394 12296 13806
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10796 6322 10824 6666
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 11164 5778 11192 6734
rect 11532 6322 11560 6734
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11716 6390 11744 6598
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11348 5778 11376 6054
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10336 800 10364 3402
rect 11624 800 11652 4490
rect 11808 4146 11836 12786
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 5370 12480 6190
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13556 4690 13584 4966
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 13372 4282 13400 4490
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 14476 3534 14504 17070
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14936 13394 14964 13670
rect 15120 13394 15148 14214
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 15488 800 15516 13330
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18064 800 18092 3470
rect 19352 800 19380 30058
rect 19996 29850 20024 30126
rect 26240 30116 26292 30122
rect 26240 30058 26292 30064
rect 25504 30048 25556 30054
rect 25504 29990 25556 29996
rect 25688 30048 25740 30054
rect 25688 29990 25740 29996
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 23480 29844 23532 29850
rect 23480 29786 23532 29792
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 23492 28966 23520 29786
rect 25516 29714 25544 29990
rect 25700 29714 25728 29990
rect 26056 29776 26108 29782
rect 26056 29718 26108 29724
rect 25504 29708 25556 29714
rect 25504 29650 25556 29656
rect 25688 29708 25740 29714
rect 25688 29650 25740 29656
rect 26068 29578 26096 29718
rect 26056 29572 26108 29578
rect 26056 29514 26108 29520
rect 23480 28960 23532 28966
rect 23480 28902 23532 28908
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 23020 24608 23072 24614
rect 23020 24550 23072 24556
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 23032 23730 23060 24550
rect 23216 23798 23244 24550
rect 23204 23792 23256 23798
rect 23204 23734 23256 23740
rect 23020 23724 23072 23730
rect 23020 23666 23072 23672
rect 24676 23656 24728 23662
rect 24676 23598 24728 23604
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 24136 18290 24164 18702
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 24320 18358 24348 18566
rect 24308 18352 24360 18358
rect 24308 18294 24360 18300
rect 24124 18284 24176 18290
rect 24124 18226 24176 18232
rect 24124 18148 24176 18154
rect 24124 18090 24176 18096
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 23112 15496 23164 15502
rect 23112 15438 23164 15444
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 23124 15026 23152 15438
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23768 15094 23796 15302
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 23112 15020 23164 15026
rect 23112 14962 23164 14968
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 20732 8294 20760 11222
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 24136 3534 24164 18090
rect 24400 11552 24452 11558
rect 24400 11494 24452 11500
rect 24412 11218 24440 11494
rect 24400 11212 24452 11218
rect 24400 11154 24452 11160
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 24596 10810 24624 11018
rect 24584 10804 24636 10810
rect 24584 10746 24636 10752
rect 24492 3596 24544 3602
rect 24492 3538 24544 3544
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 24504 800 24532 3538
rect 24688 3466 24716 23598
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 24780 18766 24808 21966
rect 26160 21486 26188 21966
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 26252 16574 26280 30058
rect 27528 30048 27580 30054
rect 27528 29990 27580 29996
rect 27540 29170 27568 29990
rect 27816 29714 27844 30194
rect 28356 30184 28408 30190
rect 28356 30126 28408 30132
rect 28368 29850 28396 30126
rect 28356 29844 28408 29850
rect 28356 29786 28408 29792
rect 32784 29782 32812 36042
rect 32876 30802 32904 38286
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34152 36780 34204 36786
rect 34152 36722 34204 36728
rect 32956 36372 33008 36378
rect 32956 36314 33008 36320
rect 32968 36106 32996 36314
rect 34164 36174 34192 36722
rect 34704 36712 34756 36718
rect 34704 36654 34756 36660
rect 34428 36576 34480 36582
rect 34428 36518 34480 36524
rect 33784 36168 33836 36174
rect 33784 36110 33836 36116
rect 34152 36168 34204 36174
rect 34152 36110 34204 36116
rect 32956 36100 33008 36106
rect 32956 36042 33008 36048
rect 32864 30796 32916 30802
rect 32864 30738 32916 30744
rect 33600 30728 33652 30734
rect 33600 30670 33652 30676
rect 32772 29776 32824 29782
rect 32772 29718 32824 29724
rect 27804 29708 27856 29714
rect 27804 29650 27856 29656
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27712 29096 27764 29102
rect 27712 29038 27764 29044
rect 30748 29096 30800 29102
rect 30748 29038 30800 29044
rect 27724 28762 27752 29038
rect 28080 29028 28132 29034
rect 28080 28970 28132 28976
rect 27712 28756 27764 28762
rect 27712 28698 27764 28704
rect 26884 26376 26936 26382
rect 26884 26318 26936 26324
rect 26896 25430 26924 26318
rect 28092 26234 28120 28970
rect 30760 28558 30788 29038
rect 33612 28558 33640 30670
rect 33796 29170 33824 36110
rect 34440 31346 34468 36518
rect 34612 35624 34664 35630
rect 34612 35566 34664 35572
rect 34428 31340 34480 31346
rect 34428 31282 34480 31288
rect 34440 30734 34468 31282
rect 34428 30728 34480 30734
rect 34428 30670 34480 30676
rect 33784 29164 33836 29170
rect 33784 29106 33836 29112
rect 33796 29050 33824 29106
rect 33704 29022 33824 29050
rect 30748 28552 30800 28558
rect 30748 28494 30800 28500
rect 33600 28552 33652 28558
rect 33600 28494 33652 28500
rect 27908 26206 28120 26234
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 26884 25424 26936 25430
rect 26884 25366 26936 25372
rect 27172 24954 27200 25842
rect 27528 25696 27580 25702
rect 27528 25638 27580 25644
rect 27540 25362 27568 25638
rect 27528 25356 27580 25362
rect 27528 25298 27580 25304
rect 27160 24948 27212 24954
rect 27160 24890 27212 24896
rect 26608 22092 26660 22098
rect 26608 22034 26660 22040
rect 26620 21690 26648 22034
rect 26608 21684 26660 21690
rect 26608 21626 26660 21632
rect 27172 20942 27200 24890
rect 27160 20936 27212 20942
rect 27160 20878 27212 20884
rect 27908 19378 27936 26206
rect 28172 25288 28224 25294
rect 28172 25230 28224 25236
rect 28184 24818 28212 25230
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 28000 24614 28028 24754
rect 28540 24744 28592 24750
rect 28540 24686 28592 24692
rect 27988 24608 28040 24614
rect 27988 24550 28040 24556
rect 28552 24410 28580 24686
rect 28540 24404 28592 24410
rect 28540 24346 28592 24352
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 26252 16546 26648 16574
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24872 10062 24900 10610
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24676 3460 24728 3466
rect 24676 3402 24728 3408
rect 7300 734 7604 762
rect 7718 0 7830 800
rect 9006 0 9118 800
rect 10294 0 10406 800
rect 11582 0 11694 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 15446 0 15558 800
rect 16734 0 16846 800
rect 18022 0 18134 800
rect 19310 0 19422 800
rect 20598 0 20710 800
rect 21886 0 21998 800
rect 23174 0 23286 800
rect 24462 0 24574 800
rect 25750 0 25862 800
rect 26620 762 26648 16546
rect 27908 15502 27936 19314
rect 27988 19168 28040 19174
rect 27988 19110 28040 19116
rect 29000 19168 29052 19174
rect 29000 19110 29052 19116
rect 28000 18834 28028 19110
rect 29012 18834 29040 19110
rect 27988 18828 28040 18834
rect 27988 18770 28040 18776
rect 29000 18828 29052 18834
rect 29000 18770 29052 18776
rect 27896 15496 27948 15502
rect 27896 15438 27948 15444
rect 30760 13938 30788 28494
rect 32128 25356 32180 25362
rect 32128 25298 32180 25304
rect 32140 24818 32168 25298
rect 32312 25152 32364 25158
rect 32312 25094 32364 25100
rect 32324 24886 32352 25094
rect 33704 24954 33732 29022
rect 33784 26920 33836 26926
rect 33784 26862 33836 26868
rect 33796 26586 33824 26862
rect 33784 26580 33836 26586
rect 33784 26522 33836 26528
rect 34624 26234 34652 35566
rect 34716 27606 34744 36654
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35360 35630 35388 49778
rect 35452 36718 35480 55694
rect 35532 45960 35584 45966
rect 35532 45902 35584 45908
rect 35440 36712 35492 36718
rect 35440 36654 35492 36660
rect 35440 36032 35492 36038
rect 35440 35974 35492 35980
rect 35348 35624 35400 35630
rect 35348 35566 35400 35572
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 35360 34610 35388 35566
rect 34796 34604 34848 34610
rect 34796 34546 34848 34552
rect 35348 34604 35400 34610
rect 35348 34546 35400 34552
rect 34704 27600 34756 27606
rect 34704 27542 34756 27548
rect 34808 27418 34836 34546
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 35452 29306 35480 35974
rect 35544 34066 35572 45902
rect 35728 45554 35756 58534
rect 35820 57390 35848 68462
rect 36096 64874 36124 71200
rect 36096 64846 37228 64874
rect 37200 59090 37228 64846
rect 37280 62280 37332 62286
rect 37280 62222 37332 62228
rect 37292 61810 37320 62222
rect 37280 61804 37332 61810
rect 37280 61746 37332 61752
rect 37384 61674 37412 71200
rect 39212 66292 39264 66298
rect 39212 66234 39264 66240
rect 37372 61668 37424 61674
rect 37372 61610 37424 61616
rect 37188 59084 37240 59090
rect 37188 59026 37240 59032
rect 38108 58404 38160 58410
rect 38108 58346 38160 58352
rect 37924 58336 37976 58342
rect 37924 58278 37976 58284
rect 37936 58002 37964 58278
rect 37924 57996 37976 58002
rect 37924 57938 37976 57944
rect 38120 57934 38148 58346
rect 38108 57928 38160 57934
rect 38108 57870 38160 57876
rect 35808 57384 35860 57390
rect 35808 57326 35860 57332
rect 38016 54664 38068 54670
rect 38016 54606 38068 54612
rect 37924 51264 37976 51270
rect 37924 51206 37976 51212
rect 35636 45526 35756 45554
rect 35636 36854 35664 45526
rect 37372 37664 37424 37670
rect 37372 37606 37424 37612
rect 37384 37330 37412 37606
rect 37372 37324 37424 37330
rect 37372 37266 37424 37272
rect 36544 37188 36596 37194
rect 36544 37130 36596 37136
rect 36636 37188 36688 37194
rect 36636 37130 36688 37136
rect 35624 36848 35676 36854
rect 35624 36790 35676 36796
rect 35532 34060 35584 34066
rect 35532 34002 35584 34008
rect 35440 29300 35492 29306
rect 35440 29242 35492 29248
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 35348 27600 35400 27606
rect 35348 27542 35400 27548
rect 34716 27390 34836 27418
rect 34716 26466 34744 27390
rect 34796 26920 34848 26926
rect 34796 26862 34848 26868
rect 34808 26586 34836 26862
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34796 26580 34848 26586
rect 34796 26522 34848 26528
rect 34716 26438 34836 26466
rect 34624 26206 34744 26234
rect 33692 24948 33744 24954
rect 33692 24890 33744 24896
rect 32312 24880 32364 24886
rect 32312 24822 32364 24828
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 31760 24676 31812 24682
rect 31760 24618 31812 24624
rect 30748 13932 30800 13938
rect 30748 13874 30800 13880
rect 30288 13252 30340 13258
rect 30288 13194 30340 13200
rect 30300 12986 30328 13194
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 27528 11144 27580 11150
rect 27528 11086 27580 11092
rect 27540 10674 27568 11086
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27896 10600 27948 10606
rect 27896 10542 27948 10548
rect 29368 10600 29420 10606
rect 29368 10542 29420 10548
rect 27908 10266 27936 10542
rect 27896 10260 27948 10266
rect 27896 10202 27948 10208
rect 29000 4752 29052 4758
rect 29000 4694 29052 4700
rect 29012 4146 29040 4694
rect 28816 4140 28868 4146
rect 28816 4082 28868 4088
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 28828 3534 28856 4082
rect 29380 3602 29408 10542
rect 29552 4616 29604 4622
rect 29552 4558 29604 4564
rect 29564 3602 29592 4558
rect 29644 4072 29696 4078
rect 29644 4014 29696 4020
rect 29368 3596 29420 3602
rect 29368 3538 29420 3544
rect 29552 3596 29604 3602
rect 29552 3538 29604 3544
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 26896 870 27108 898
rect 26896 762 26924 870
rect 27080 800 27108 870
rect 29656 800 29684 4014
rect 26620 734 26924 762
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 29614 0 29726 800
rect 30902 0 31014 800
rect 31772 762 31800 24618
rect 33704 17678 33732 24890
rect 34716 19378 34744 26206
rect 34808 24206 34836 26438
rect 35360 26382 35388 27542
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34796 24200 34848 24206
rect 34796 24142 34848 24148
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 35360 22642 35388 26318
rect 35452 24614 35480 29242
rect 35544 27470 35572 34002
rect 35636 29646 35664 36790
rect 36084 36780 36136 36786
rect 36084 36722 36136 36728
rect 36096 36174 36124 36722
rect 36556 36174 36584 37130
rect 36648 36922 36676 37130
rect 37372 37120 37424 37126
rect 37372 37062 37424 37068
rect 36636 36916 36688 36922
rect 36636 36858 36688 36864
rect 37384 36786 37412 37062
rect 37936 36854 37964 51206
rect 38028 36854 38056 54606
rect 38200 42220 38252 42226
rect 38200 42162 38252 42168
rect 37648 36848 37700 36854
rect 37648 36790 37700 36796
rect 37924 36848 37976 36854
rect 37924 36790 37976 36796
rect 38016 36848 38068 36854
rect 38016 36790 38068 36796
rect 37372 36780 37424 36786
rect 37372 36722 37424 36728
rect 37384 36174 37412 36722
rect 36084 36168 36136 36174
rect 36084 36110 36136 36116
rect 36544 36168 36596 36174
rect 36544 36110 36596 36116
rect 37372 36168 37424 36174
rect 37372 36110 37424 36116
rect 35900 36032 35952 36038
rect 35900 35974 35952 35980
rect 35912 35698 35940 35974
rect 35900 35692 35952 35698
rect 35900 35634 35952 35640
rect 35912 34610 35940 35634
rect 37384 34610 37412 36110
rect 35900 34604 35952 34610
rect 35900 34546 35952 34552
rect 37372 34604 37424 34610
rect 37372 34546 37424 34552
rect 35912 33998 35940 34546
rect 36452 34060 36504 34066
rect 36452 34002 36504 34008
rect 35900 33992 35952 33998
rect 35900 33934 35952 33940
rect 35624 29640 35676 29646
rect 35624 29582 35676 29588
rect 35532 27464 35584 27470
rect 35532 27406 35584 27412
rect 35440 24608 35492 24614
rect 35440 24550 35492 24556
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35544 22098 35572 27406
rect 35636 26234 35664 29582
rect 35636 26206 35756 26234
rect 35728 25294 35756 26206
rect 35716 25288 35768 25294
rect 35716 25230 35768 25236
rect 35532 22092 35584 22098
rect 35532 22034 35584 22040
rect 36464 21554 36492 34002
rect 37384 33998 37412 34546
rect 37372 33992 37424 33998
rect 37372 33934 37424 33940
rect 37660 29714 37688 36790
rect 38212 34542 38240 42162
rect 38844 42152 38896 42158
rect 38844 42094 38896 42100
rect 38660 36780 38712 36786
rect 38660 36722 38712 36728
rect 38672 35894 38700 36722
rect 38580 35866 38700 35894
rect 38200 34536 38252 34542
rect 38200 34478 38252 34484
rect 37648 29708 37700 29714
rect 37648 29650 37700 29656
rect 36452 21548 36504 21554
rect 36452 21490 36504 21496
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34704 19372 34756 19378
rect 34704 19314 34756 19320
rect 35716 19236 35768 19242
rect 35716 19178 35768 19184
rect 35532 19168 35584 19174
rect 35532 19110 35584 19116
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 35544 18834 35572 19110
rect 35728 18834 35756 19178
rect 35532 18828 35584 18834
rect 35532 18770 35584 18776
rect 35716 18828 35768 18834
rect 35716 18770 35768 18776
rect 37188 18828 37240 18834
rect 37188 18770 37240 18776
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 33692 17672 33744 17678
rect 33692 17614 33744 17620
rect 36820 17672 36872 17678
rect 36820 17614 36872 17620
rect 36832 17202 36860 17614
rect 36820 17196 36872 17202
rect 36820 17138 36872 17144
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 36360 14408 36412 14414
rect 36360 14350 36412 14356
rect 35808 14272 35860 14278
rect 35808 14214 35860 14220
rect 31944 14000 31996 14006
rect 31944 13942 31996 13948
rect 31956 13394 31984 13942
rect 32128 13864 32180 13870
rect 32128 13806 32180 13812
rect 32140 13394 32168 13806
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 35820 13394 35848 14214
rect 36372 13462 36400 14350
rect 36360 13456 36412 13462
rect 36360 13398 36412 13404
rect 31944 13388 31996 13394
rect 31944 13330 31996 13336
rect 32128 13388 32180 13394
rect 32128 13330 32180 13336
rect 35808 13388 35860 13394
rect 35808 13330 35860 13336
rect 36084 13388 36136 13394
rect 36084 13330 36136 13336
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 32048 870 32260 898
rect 32048 762 32076 870
rect 32232 800 32260 870
rect 36096 800 36124 13330
rect 37200 3534 37228 18770
rect 38212 10674 38240 34478
rect 38580 31346 38608 35866
rect 38568 31340 38620 31346
rect 38568 31282 38620 31288
rect 38580 29170 38608 31282
rect 38856 31278 38884 42094
rect 39224 37262 39252 66234
rect 40144 52630 40172 71318
rect 41206 71200 41318 71318
rect 41432 71318 42606 71346
rect 40316 58540 40368 58546
rect 40316 58482 40368 58488
rect 40328 58002 40356 58482
rect 40316 57996 40368 58002
rect 40316 57938 40368 57944
rect 40132 52624 40184 52630
rect 40132 52566 40184 52572
rect 39212 37256 39264 37262
rect 39212 37198 39264 37204
rect 40328 36854 40356 57938
rect 40776 54596 40828 54602
rect 40776 54538 40828 54544
rect 40684 52896 40736 52902
rect 40684 52838 40736 52844
rect 40696 52562 40724 52838
rect 40684 52556 40736 52562
rect 40684 52498 40736 52504
rect 40788 52018 40816 54538
rect 40868 52420 40920 52426
rect 40868 52362 40920 52368
rect 40880 52154 40908 52362
rect 40868 52148 40920 52154
rect 40868 52090 40920 52096
rect 40776 52012 40828 52018
rect 40776 51954 40828 51960
rect 40788 46986 40816 51954
rect 40776 46980 40828 46986
rect 40776 46922 40828 46928
rect 40788 45554 40816 46922
rect 41432 46510 41460 71318
rect 42494 71200 42606 71318
rect 43782 71200 43894 72000
rect 45070 71200 45182 72000
rect 46358 71346 46470 72000
rect 45572 71318 46470 71346
rect 43352 63368 43404 63374
rect 43352 63310 43404 63316
rect 43628 63368 43680 63374
rect 43628 63310 43680 63316
rect 43364 62898 43392 63310
rect 43640 62898 43668 63310
rect 43812 63232 43864 63238
rect 43812 63174 43864 63180
rect 43824 62966 43852 63174
rect 43812 62960 43864 62966
rect 43812 62902 43864 62908
rect 43352 62892 43404 62898
rect 43352 62834 43404 62840
rect 43628 62892 43680 62898
rect 43628 62834 43680 62840
rect 41420 46504 41472 46510
rect 41420 46446 41472 46452
rect 42432 46504 42484 46510
rect 42432 46446 42484 46452
rect 41972 46368 42024 46374
rect 41972 46310 42024 46316
rect 41984 46034 42012 46310
rect 42444 46034 42472 46446
rect 41972 46028 42024 46034
rect 41972 45970 42024 45976
rect 42432 46028 42484 46034
rect 42432 45970 42484 45976
rect 40696 45526 40816 45554
rect 40316 36848 40368 36854
rect 40316 36790 40368 36796
rect 40328 32910 40356 36790
rect 40696 35766 40724 45526
rect 43364 36378 43392 62834
rect 45572 61334 45600 71318
rect 46358 71200 46470 71318
rect 47646 71200 47758 72000
rect 48934 71200 49046 72000
rect 50222 71346 50334 72000
rect 49896 71318 50334 71346
rect 49424 68196 49476 68202
rect 49424 68138 49476 68144
rect 46848 68128 46900 68134
rect 46848 68070 46900 68076
rect 45836 61600 45888 61606
rect 45836 61542 45888 61548
rect 45560 61328 45612 61334
rect 45560 61270 45612 61276
rect 45848 61266 45876 61542
rect 45836 61260 45888 61266
rect 45836 61202 45888 61208
rect 46020 61124 46072 61130
rect 46020 61066 46072 61072
rect 46032 60858 46060 61066
rect 46020 60852 46072 60858
rect 46020 60794 46072 60800
rect 45928 60716 45980 60722
rect 45928 60658 45980 60664
rect 45940 59634 45968 60658
rect 45928 59628 45980 59634
rect 45928 59570 45980 59576
rect 43444 50924 43496 50930
rect 43444 50866 43496 50872
rect 43352 36372 43404 36378
rect 43352 36314 43404 36320
rect 40684 35760 40736 35766
rect 40684 35702 40736 35708
rect 41420 35692 41472 35698
rect 41420 35634 41472 35640
rect 41432 34066 41460 35634
rect 43260 34604 43312 34610
rect 43260 34546 43312 34552
rect 41420 34060 41472 34066
rect 41420 34002 41472 34008
rect 40316 32904 40368 32910
rect 40316 32846 40368 32852
rect 38844 31272 38896 31278
rect 38844 31214 38896 31220
rect 38660 29300 38712 29306
rect 38660 29242 38712 29248
rect 38568 29164 38620 29170
rect 38568 29106 38620 29112
rect 38672 29034 38700 29242
rect 38660 29028 38712 29034
rect 38660 28970 38712 28976
rect 38476 17740 38528 17746
rect 38476 17682 38528 17688
rect 38200 10668 38252 10674
rect 38200 10610 38252 10616
rect 38212 10062 38240 10610
rect 38292 10464 38344 10470
rect 38292 10406 38344 10412
rect 38200 10056 38252 10062
rect 38200 9998 38252 10004
rect 38304 9654 38332 10406
rect 38292 9648 38344 9654
rect 38292 9590 38344 9596
rect 38488 6914 38516 17682
rect 38856 14482 38884 31214
rect 40132 28484 40184 28490
rect 40132 28426 40184 28432
rect 38844 14476 38896 14482
rect 38844 14418 38896 14424
rect 40040 12232 40092 12238
rect 40040 12174 40092 12180
rect 40052 11762 40080 12174
rect 40040 11756 40092 11762
rect 40040 11698 40092 11704
rect 40144 11150 40172 28426
rect 41432 26234 41460 34002
rect 42432 33448 42484 33454
rect 42432 33390 42484 33396
rect 42444 33114 42472 33390
rect 42432 33108 42484 33114
rect 42432 33050 42484 33056
rect 41432 26206 41552 26234
rect 41524 12238 41552 26206
rect 41512 12232 41564 12238
rect 41512 12174 41564 12180
rect 41880 12096 41932 12102
rect 41880 12038 41932 12044
rect 40224 11688 40276 11694
rect 40224 11630 40276 11636
rect 40236 11354 40264 11630
rect 41696 11552 41748 11558
rect 41696 11494 41748 11500
rect 40224 11348 40276 11354
rect 40224 11290 40276 11296
rect 41708 11218 41736 11494
rect 41892 11218 41920 12038
rect 41696 11212 41748 11218
rect 41696 11154 41748 11160
rect 41880 11212 41932 11218
rect 41880 11154 41932 11160
rect 40132 11144 40184 11150
rect 40132 11086 40184 11092
rect 40144 10674 40172 11086
rect 40132 10668 40184 10674
rect 40132 10610 40184 10616
rect 38844 10464 38896 10470
rect 38844 10406 38896 10412
rect 38660 9512 38712 9518
rect 38660 9454 38712 9460
rect 37384 6886 38516 6914
rect 37188 3528 37240 3534
rect 37188 3470 37240 3476
rect 37384 800 37412 6886
rect 38672 800 38700 9454
rect 38856 9450 38884 10406
rect 38844 9444 38896 9450
rect 38844 9386 38896 9392
rect 43272 6866 43300 34546
rect 43364 33590 43392 36314
rect 43456 36242 43484 50866
rect 44916 47048 44968 47054
rect 44916 46990 44968 46996
rect 44928 42226 44956 46990
rect 45008 43104 45060 43110
rect 45008 43046 45060 43052
rect 45020 42770 45048 43046
rect 46860 42770 46888 68070
rect 48964 67924 49016 67930
rect 48964 67866 49016 67872
rect 48976 62830 49004 67866
rect 48964 62824 49016 62830
rect 48964 62766 49016 62772
rect 49240 56840 49292 56846
rect 49240 56782 49292 56788
rect 49252 56370 49280 56782
rect 49240 56364 49292 56370
rect 49240 56306 49292 56312
rect 49240 56228 49292 56234
rect 49240 56170 49292 56176
rect 49252 55962 49280 56170
rect 49240 55956 49292 55962
rect 49240 55898 49292 55904
rect 48688 55752 48740 55758
rect 48688 55694 48740 55700
rect 48700 55282 48728 55694
rect 48688 55276 48740 55282
rect 48688 55218 48740 55224
rect 48872 55208 48924 55214
rect 48872 55150 48924 55156
rect 48884 54874 48912 55150
rect 48872 54868 48924 54874
rect 48872 54810 48924 54816
rect 48596 54664 48648 54670
rect 48596 54606 48648 54612
rect 48608 51270 48636 54606
rect 48596 51264 48648 51270
rect 48596 51206 48648 51212
rect 48964 51264 49016 51270
rect 48964 51206 49016 51212
rect 47768 47592 47820 47598
rect 47768 47534 47820 47540
rect 47780 47258 47808 47534
rect 47768 47252 47820 47258
rect 47768 47194 47820 47200
rect 45008 42764 45060 42770
rect 45008 42706 45060 42712
rect 46848 42764 46900 42770
rect 46848 42706 46900 42712
rect 48976 42702 49004 51206
rect 49436 47734 49464 68138
rect 49896 67930 49924 71318
rect 50222 71200 50334 71318
rect 51510 71200 51622 72000
rect 52798 71200 52910 72000
rect 54086 71200 54198 72000
rect 55374 71200 55486 72000
rect 56662 71200 56774 72000
rect 57950 71200 58062 72000
rect 59238 71200 59350 72000
rect 60526 71200 60638 72000
rect 61814 71200 61926 72000
rect 63102 71200 63214 72000
rect 64390 71346 64502 72000
rect 65678 71346 65790 72000
rect 63604 71318 64502 71346
rect 50294 69660 50602 69680
rect 50294 69658 50300 69660
rect 50356 69658 50380 69660
rect 50436 69658 50460 69660
rect 50516 69658 50540 69660
rect 50596 69658 50602 69660
rect 50356 69606 50358 69658
rect 50538 69606 50540 69658
rect 50294 69604 50300 69606
rect 50356 69604 50380 69606
rect 50436 69604 50460 69606
rect 50516 69604 50540 69606
rect 50596 69604 50602 69606
rect 50294 69584 50602 69604
rect 50294 68572 50602 68592
rect 50294 68570 50300 68572
rect 50356 68570 50380 68572
rect 50436 68570 50460 68572
rect 50516 68570 50540 68572
rect 50596 68570 50602 68572
rect 50356 68518 50358 68570
rect 50538 68518 50540 68570
rect 50294 68516 50300 68518
rect 50356 68516 50380 68518
rect 50436 68516 50460 68518
rect 50516 68516 50540 68518
rect 50596 68516 50602 68518
rect 50294 68496 50602 68516
rect 50620 68332 50672 68338
rect 50620 68274 50672 68280
rect 49884 67924 49936 67930
rect 49884 67866 49936 67872
rect 50294 67484 50602 67504
rect 50294 67482 50300 67484
rect 50356 67482 50380 67484
rect 50436 67482 50460 67484
rect 50516 67482 50540 67484
rect 50596 67482 50602 67484
rect 50356 67430 50358 67482
rect 50538 67430 50540 67482
rect 50294 67428 50300 67430
rect 50356 67428 50380 67430
rect 50436 67428 50460 67430
rect 50516 67428 50540 67430
rect 50596 67428 50602 67430
rect 50294 67408 50602 67428
rect 50294 66396 50602 66416
rect 50294 66394 50300 66396
rect 50356 66394 50380 66396
rect 50436 66394 50460 66396
rect 50516 66394 50540 66396
rect 50596 66394 50602 66396
rect 50356 66342 50358 66394
rect 50538 66342 50540 66394
rect 50294 66340 50300 66342
rect 50356 66340 50380 66342
rect 50436 66340 50460 66342
rect 50516 66340 50540 66342
rect 50596 66340 50602 66342
rect 50294 66320 50602 66340
rect 50294 65308 50602 65328
rect 50294 65306 50300 65308
rect 50356 65306 50380 65308
rect 50436 65306 50460 65308
rect 50516 65306 50540 65308
rect 50596 65306 50602 65308
rect 50356 65254 50358 65306
rect 50538 65254 50540 65306
rect 50294 65252 50300 65254
rect 50356 65252 50380 65254
rect 50436 65252 50460 65254
rect 50516 65252 50540 65254
rect 50596 65252 50602 65254
rect 50294 65232 50602 65252
rect 50294 64220 50602 64240
rect 50294 64218 50300 64220
rect 50356 64218 50380 64220
rect 50436 64218 50460 64220
rect 50516 64218 50540 64220
rect 50596 64218 50602 64220
rect 50356 64166 50358 64218
rect 50538 64166 50540 64218
rect 50294 64164 50300 64166
rect 50356 64164 50380 64166
rect 50436 64164 50460 64166
rect 50516 64164 50540 64166
rect 50596 64164 50602 64166
rect 50294 64144 50602 64164
rect 50294 63132 50602 63152
rect 50294 63130 50300 63132
rect 50356 63130 50380 63132
rect 50436 63130 50460 63132
rect 50516 63130 50540 63132
rect 50596 63130 50602 63132
rect 50356 63078 50358 63130
rect 50538 63078 50540 63130
rect 50294 63076 50300 63078
rect 50356 63076 50380 63078
rect 50436 63076 50460 63078
rect 50516 63076 50540 63078
rect 50596 63076 50602 63078
rect 50294 63056 50602 63076
rect 50294 62044 50602 62064
rect 50294 62042 50300 62044
rect 50356 62042 50380 62044
rect 50436 62042 50460 62044
rect 50516 62042 50540 62044
rect 50596 62042 50602 62044
rect 50356 61990 50358 62042
rect 50538 61990 50540 62042
rect 50294 61988 50300 61990
rect 50356 61988 50380 61990
rect 50436 61988 50460 61990
rect 50516 61988 50540 61990
rect 50596 61988 50602 61990
rect 50294 61968 50602 61988
rect 50294 60956 50602 60976
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60880 50602 60900
rect 50294 59868 50602 59888
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59792 50602 59812
rect 50294 58780 50602 58800
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58704 50602 58724
rect 50294 57692 50602 57712
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57616 50602 57636
rect 50294 56604 50602 56624
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56528 50602 56548
rect 50294 55516 50602 55536
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55440 50602 55460
rect 50632 55350 50660 68274
rect 51552 68134 51580 71200
rect 52828 69012 52880 69018
rect 52828 68954 52880 68960
rect 51540 68128 51592 68134
rect 51540 68070 51592 68076
rect 50620 55344 50672 55350
rect 50620 55286 50672 55292
rect 50294 54428 50602 54448
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54352 50602 54372
rect 50294 53340 50602 53360
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53264 50602 53284
rect 50294 52252 50602 52272
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52176 50602 52196
rect 50988 51808 51040 51814
rect 50988 51750 51040 51756
rect 51000 51474 51028 51750
rect 52840 51474 52868 68954
rect 54128 68202 54156 71200
rect 56704 69018 56732 71200
rect 56692 69012 56744 69018
rect 56692 68954 56744 68960
rect 54116 68196 54168 68202
rect 54116 68138 54168 68144
rect 57992 64874 58020 71200
rect 62764 69216 62816 69222
rect 62764 69158 62816 69164
rect 62028 68808 62080 68814
rect 62028 68750 62080 68756
rect 57992 64846 59124 64874
rect 54116 61872 54168 61878
rect 54116 61814 54168 61820
rect 54128 61198 54156 61814
rect 55312 61600 55364 61606
rect 55312 61542 55364 61548
rect 55324 61266 55352 61542
rect 55312 61260 55364 61266
rect 55312 61202 55364 61208
rect 54116 61192 54168 61198
rect 54116 61134 54168 61140
rect 54852 60104 54904 60110
rect 54852 60046 54904 60052
rect 54864 59634 54892 60046
rect 54852 59628 54904 59634
rect 54852 59570 54904 59576
rect 50988 51468 51040 51474
rect 50988 51410 51040 51416
rect 52828 51468 52880 51474
rect 52828 51410 52880 51416
rect 51172 51332 51224 51338
rect 51172 51274 51224 51280
rect 50294 51164 50602 51184
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51088 50602 51108
rect 51184 51066 51212 51274
rect 51172 51060 51224 51066
rect 51172 51002 51224 51008
rect 50294 50076 50602 50096
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50000 50602 50020
rect 54116 49224 54168 49230
rect 54116 49166 54168 49172
rect 50294 48988 50602 49008
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48912 50602 48932
rect 54128 48754 54156 49166
rect 51080 48748 51132 48754
rect 51080 48690 51132 48696
rect 54116 48748 54168 48754
rect 54116 48690 54168 48696
rect 50294 47900 50602 47920
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47824 50602 47844
rect 49424 47728 49476 47734
rect 49424 47670 49476 47676
rect 50294 46812 50602 46832
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46736 50602 46756
rect 51092 46102 51120 48690
rect 58072 47116 58124 47122
rect 58072 47058 58124 47064
rect 56508 47048 56560 47054
rect 56508 46990 56560 46996
rect 51080 46096 51132 46102
rect 51080 46038 51132 46044
rect 50294 45724 50602 45744
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45648 50602 45668
rect 50294 44636 50602 44656
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44560 50602 44580
rect 50294 43548 50602 43568
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43472 50602 43492
rect 52736 43104 52788 43110
rect 52736 43046 52788 43052
rect 52748 42770 52776 43046
rect 52736 42764 52788 42770
rect 52736 42706 52788 42712
rect 48964 42696 49016 42702
rect 48964 42638 49016 42644
rect 45008 42628 45060 42634
rect 45008 42570 45060 42576
rect 45020 42362 45048 42570
rect 50294 42460 50602 42480
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42384 50602 42404
rect 45008 42356 45060 42362
rect 45008 42298 45060 42304
rect 44916 42220 44968 42226
rect 44916 42162 44968 42168
rect 50294 41372 50602 41392
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41296 50602 41316
rect 50294 40284 50602 40304
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40208 50602 40228
rect 50294 39196 50602 39216
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39120 50602 39140
rect 50294 38108 50602 38128
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38032 50602 38052
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 43444 36236 43496 36242
rect 43444 36178 43496 36184
rect 43352 33584 43404 33590
rect 43352 33526 43404 33532
rect 43456 32434 43484 36178
rect 45192 36168 45244 36174
rect 45192 36110 45244 36116
rect 45204 35698 45232 36110
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 45192 35692 45244 35698
rect 45192 35634 45244 35640
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 49148 33992 49200 33998
rect 49148 33934 49200 33940
rect 55496 33992 55548 33998
rect 55496 33934 55548 33940
rect 49160 33522 49188 33934
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 55508 33522 55536 33934
rect 49148 33516 49200 33522
rect 49148 33458 49200 33464
rect 55496 33516 55548 33522
rect 55496 33458 55548 33464
rect 49332 33448 49384 33454
rect 49332 33390 49384 33396
rect 55680 33448 55732 33454
rect 55680 33390 55732 33396
rect 49344 33114 49372 33390
rect 55692 33114 55720 33390
rect 49332 33108 49384 33114
rect 49332 33050 49384 33056
rect 55680 33108 55732 33114
rect 55680 33050 55732 33056
rect 49056 32904 49108 32910
rect 49056 32846 49108 32852
rect 49068 32570 49096 32846
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 49056 32564 49108 32570
rect 49056 32506 49108 32512
rect 43444 32428 43496 32434
rect 43444 32370 43496 32376
rect 44548 32360 44600 32366
rect 44548 32302 44600 32308
rect 44180 32292 44232 32298
rect 44180 32234 44232 32240
rect 44192 16574 44220 32234
rect 44560 32026 44588 32302
rect 44548 32020 44600 32026
rect 44548 31962 44600 31968
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 51080 30048 51132 30054
rect 51080 29990 51132 29996
rect 50988 29640 51040 29646
rect 50988 29582 51040 29588
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 51000 29034 51028 29582
rect 50988 29028 51040 29034
rect 50988 28970 51040 28976
rect 51092 28626 51120 29990
rect 51724 29572 51776 29578
rect 51724 29514 51776 29520
rect 53380 29572 53432 29578
rect 53380 29514 53432 29520
rect 51264 29504 51316 29510
rect 51264 29446 51316 29452
rect 51276 28626 51304 29446
rect 51736 29238 51764 29514
rect 51724 29232 51776 29238
rect 51724 29174 51776 29180
rect 51080 28620 51132 28626
rect 51080 28562 51132 28568
rect 51264 28620 51316 28626
rect 51264 28562 51316 28568
rect 52920 28484 52972 28490
rect 52920 28426 52972 28432
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 50528 28008 50580 28014
rect 50528 27950 50580 27956
rect 50540 27674 50568 27950
rect 50528 27668 50580 27674
rect 50528 27610 50580 27616
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 52184 22568 52236 22574
rect 52184 22510 52236 22516
rect 52196 22234 52224 22510
rect 52184 22228 52236 22234
rect 52184 22170 52236 22176
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 52932 17882 52960 28426
rect 53392 19310 53420 29514
rect 55772 26784 55824 26790
rect 55772 26726 55824 26732
rect 55784 26450 55812 26726
rect 55772 26444 55824 26450
rect 55772 26386 55824 26392
rect 55956 26308 56008 26314
rect 55956 26250 56008 26256
rect 55968 26042 55996 26250
rect 55956 26036 56008 26042
rect 55956 25978 56008 25984
rect 56520 25906 56548 46990
rect 58084 46578 58112 47058
rect 58072 46572 58124 46578
rect 58072 46514 58124 46520
rect 57428 42016 57480 42022
rect 57428 41958 57480 41964
rect 57440 41682 57468 41958
rect 59096 41682 59124 64846
rect 61936 47456 61988 47462
rect 61936 47398 61988 47404
rect 61948 47122 61976 47398
rect 61936 47116 61988 47122
rect 61936 47058 61988 47064
rect 60924 46572 60976 46578
rect 60924 46514 60976 46520
rect 60832 45416 60884 45422
rect 60832 45358 60884 45364
rect 60844 45082 60872 45358
rect 60832 45076 60884 45082
rect 60832 45018 60884 45024
rect 60556 44872 60608 44878
rect 60556 44814 60608 44820
rect 60280 43784 60332 43790
rect 60280 43726 60332 43732
rect 60292 43314 60320 43726
rect 60280 43308 60332 43314
rect 60280 43250 60332 43256
rect 60464 43240 60516 43246
rect 60464 43182 60516 43188
rect 60476 42906 60504 43182
rect 60464 42900 60516 42906
rect 60464 42842 60516 42848
rect 60568 42702 60596 44814
rect 59728 42696 59780 42702
rect 59728 42638 59780 42644
rect 60556 42696 60608 42702
rect 60556 42638 60608 42644
rect 57428 41676 57480 41682
rect 57428 41618 57480 41624
rect 59084 41676 59136 41682
rect 59084 41618 59136 41624
rect 56784 41608 56836 41614
rect 56784 41550 56836 41556
rect 56796 31278 56824 41550
rect 57336 33448 57388 33454
rect 57336 33390 57388 33396
rect 56784 31272 56836 31278
rect 56784 31214 56836 31220
rect 56508 25900 56560 25906
rect 56508 25842 56560 25848
rect 54576 22568 54628 22574
rect 54576 22510 54628 22516
rect 53380 19304 53432 19310
rect 53380 19246 53432 19252
rect 52920 17876 52972 17882
rect 52920 17818 52972 17824
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 44192 16546 44680 16574
rect 44088 10464 44140 10470
rect 44088 10406 44140 10412
rect 44100 10198 44128 10406
rect 44088 10192 44140 10198
rect 44088 10134 44140 10140
rect 43260 6860 43312 6866
rect 43260 6802 43312 6808
rect 43272 6322 43300 6802
rect 43260 6316 43312 6322
rect 43260 6258 43312 6264
rect 43628 6112 43680 6118
rect 43628 6054 43680 6060
rect 43444 5704 43496 5710
rect 43444 5646 43496 5652
rect 43456 5234 43484 5646
rect 43640 5302 43668 6054
rect 43628 5296 43680 5302
rect 43628 5238 43680 5244
rect 43444 5228 43496 5234
rect 43444 5170 43496 5176
rect 31772 734 32076 762
rect 32190 0 32302 800
rect 33478 0 33590 800
rect 34766 0 34878 800
rect 36054 0 36166 800
rect 37342 0 37454 800
rect 38630 0 38742 800
rect 39918 0 40030 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43782 0 43894 800
rect 44652 762 44680 16546
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 45008 10464 45060 10470
rect 45008 10406 45060 10412
rect 45020 10130 45048 10406
rect 45008 10124 45060 10130
rect 45008 10066 45060 10072
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 47768 8288 47820 8294
rect 47768 8230 47820 8236
rect 47780 7954 47808 8230
rect 47768 7948 47820 7954
rect 47768 7890 47820 7896
rect 47124 7880 47176 7886
rect 47124 7822 47176 7828
rect 47136 6866 47164 7822
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 47124 6860 47176 6866
rect 47124 6802 47176 6808
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 54588 3670 54616 22510
rect 56324 22432 56376 22438
rect 56324 22374 56376 22380
rect 56336 22098 56364 22374
rect 56324 22092 56376 22098
rect 56324 22034 56376 22040
rect 56324 21956 56376 21962
rect 56324 21898 56376 21904
rect 56336 21690 56364 21898
rect 56324 21684 56376 21690
rect 56324 21626 56376 21632
rect 56520 21554 56548 25842
rect 56508 21548 56560 21554
rect 56508 21490 56560 21496
rect 57244 11076 57296 11082
rect 57244 11018 57296 11024
rect 54576 3664 54628 3670
rect 54576 3606 54628 3612
rect 56048 3596 56100 3602
rect 56048 3538 56100 3544
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 44928 870 45140 898
rect 44928 762 44956 870
rect 45112 800 45140 870
rect 56060 800 56088 3538
rect 57256 3482 57284 11018
rect 57348 3602 57376 33390
rect 58164 31272 58216 31278
rect 58164 31214 58216 31220
rect 58072 26784 58124 26790
rect 58072 26726 58124 26732
rect 58084 26450 58112 26726
rect 58072 26444 58124 26450
rect 58072 26386 58124 26392
rect 57612 26308 57664 26314
rect 57612 26250 57664 26256
rect 57624 3602 57652 26250
rect 58176 25906 58204 31214
rect 59740 30734 59768 42638
rect 60936 37262 60964 46514
rect 61016 45960 61068 45966
rect 61016 45902 61068 45908
rect 61028 45558 61056 45902
rect 61016 45552 61068 45558
rect 61016 45494 61068 45500
rect 62040 43246 62068 68750
rect 62776 59702 62804 69158
rect 62764 59696 62816 59702
rect 62764 59638 62816 59644
rect 63500 57928 63552 57934
rect 63500 57870 63552 57876
rect 63512 57458 63540 57870
rect 63500 57452 63552 57458
rect 63500 57394 63552 57400
rect 63604 56506 63632 71318
rect 64390 71200 64502 71318
rect 65352 71318 65790 71346
rect 65352 68814 65380 71318
rect 65678 71200 65790 71318
rect 66966 71200 67078 72000
rect 68254 71200 68366 72000
rect 69542 71200 69654 72000
rect 66074 70136 66130 70145
rect 66074 70071 66130 70080
rect 66088 69222 66116 70071
rect 66076 69216 66128 69222
rect 66076 69158 66128 69164
rect 65654 69116 65962 69136
rect 65654 69114 65660 69116
rect 65716 69114 65740 69116
rect 65796 69114 65820 69116
rect 65876 69114 65900 69116
rect 65956 69114 65962 69116
rect 65716 69062 65718 69114
rect 65898 69062 65900 69114
rect 65654 69060 65660 69062
rect 65716 69060 65740 69062
rect 65796 69060 65820 69062
rect 65876 69060 65900 69062
rect 65956 69060 65962 69062
rect 65654 69040 65962 69060
rect 65340 68808 65392 68814
rect 65340 68750 65392 68756
rect 67008 68338 67036 71200
rect 66996 68332 67048 68338
rect 66996 68274 67048 68280
rect 65654 68028 65962 68048
rect 65654 68026 65660 68028
rect 65716 68026 65740 68028
rect 65796 68026 65820 68028
rect 65876 68026 65900 68028
rect 65956 68026 65962 68028
rect 65716 67974 65718 68026
rect 65898 67974 65900 68026
rect 65654 67972 65660 67974
rect 65716 67972 65740 67974
rect 65796 67972 65820 67974
rect 65876 67972 65900 67974
rect 65956 67972 65962 67974
rect 65654 67952 65962 67972
rect 65338 67416 65394 67425
rect 65338 67351 65394 67360
rect 65352 66298 65380 67351
rect 65654 66940 65962 66960
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66864 65962 66884
rect 65340 66292 65392 66298
rect 65340 66234 65392 66240
rect 64878 66056 64934 66065
rect 64878 65991 64934 66000
rect 64892 61130 64920 65991
rect 65654 65852 65962 65872
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65776 65962 65796
rect 65654 64764 65962 64784
rect 65654 64762 65660 64764
rect 65716 64762 65740 64764
rect 65796 64762 65820 64764
rect 65876 64762 65900 64764
rect 65956 64762 65962 64764
rect 65716 64710 65718 64762
rect 65898 64710 65900 64762
rect 65654 64708 65660 64710
rect 65716 64708 65740 64710
rect 65796 64708 65820 64710
rect 65876 64708 65900 64710
rect 65956 64708 65962 64710
rect 65654 64688 65962 64708
rect 66074 64696 66130 64705
rect 66074 64631 66130 64640
rect 65654 63676 65962 63696
rect 65654 63674 65660 63676
rect 65716 63674 65740 63676
rect 65796 63674 65820 63676
rect 65876 63674 65900 63676
rect 65956 63674 65962 63676
rect 65716 63622 65718 63674
rect 65898 63622 65900 63674
rect 65654 63620 65660 63622
rect 65716 63620 65740 63622
rect 65796 63620 65820 63622
rect 65876 63620 65900 63622
rect 65956 63620 65962 63622
rect 65654 63600 65962 63620
rect 65654 62588 65962 62608
rect 65654 62586 65660 62588
rect 65716 62586 65740 62588
rect 65796 62586 65820 62588
rect 65876 62586 65900 62588
rect 65956 62586 65962 62588
rect 65716 62534 65718 62586
rect 65898 62534 65900 62586
rect 65654 62532 65660 62534
rect 65716 62532 65740 62534
rect 65796 62532 65820 62534
rect 65876 62532 65900 62534
rect 65956 62532 65962 62534
rect 65654 62512 65962 62532
rect 65430 61976 65486 61985
rect 65430 61911 65486 61920
rect 64880 61124 64932 61130
rect 64880 61066 64932 61072
rect 64512 58472 64564 58478
rect 64512 58414 64564 58420
rect 64524 58138 64552 58414
rect 64512 58132 64564 58138
rect 64512 58074 64564 58080
rect 63684 57996 63736 58002
rect 63684 57938 63736 57944
rect 63592 56500 63644 56506
rect 63592 56442 63644 56448
rect 63696 55758 63724 57938
rect 64236 57792 64288 57798
rect 64236 57734 64288 57740
rect 64248 57526 64276 57734
rect 64236 57520 64288 57526
rect 64236 57462 64288 57468
rect 63960 56840 64012 56846
rect 63960 56782 64012 56788
rect 63972 56370 64000 56782
rect 64420 56500 64472 56506
rect 64420 56442 64472 56448
rect 63960 56364 64012 56370
rect 63960 56306 64012 56312
rect 64432 56302 64460 56442
rect 64236 56296 64288 56302
rect 64236 56238 64288 56244
rect 64420 56296 64472 56302
rect 64420 56238 64472 56244
rect 64248 55962 64276 56238
rect 64236 55956 64288 55962
rect 64236 55898 64288 55904
rect 63684 55752 63736 55758
rect 63684 55694 63736 55700
rect 64696 55752 64748 55758
rect 64696 55694 64748 55700
rect 64972 55752 65024 55758
rect 64972 55694 65024 55700
rect 63592 55616 63644 55622
rect 63592 55558 63644 55564
rect 63224 55072 63276 55078
rect 63224 55014 63276 55020
rect 63236 54738 63264 55014
rect 63604 54738 63632 55558
rect 63224 54732 63276 54738
rect 63224 54674 63276 54680
rect 63592 54732 63644 54738
rect 63592 54674 63644 54680
rect 62120 46980 62172 46986
rect 62120 46922 62172 46928
rect 62132 46714 62160 46922
rect 62120 46708 62172 46714
rect 62120 46650 62172 46656
rect 62028 43240 62080 43246
rect 62028 43182 62080 43188
rect 61384 40112 61436 40118
rect 61384 40054 61436 40060
rect 60924 37256 60976 37262
rect 60924 37198 60976 37204
rect 61292 37256 61344 37262
rect 61292 37198 61344 37204
rect 61304 35630 61332 37198
rect 61396 35766 61424 40054
rect 64708 38962 64736 55694
rect 64984 55282 65012 55694
rect 65156 55616 65208 55622
rect 65156 55558 65208 55564
rect 65168 55350 65196 55558
rect 65156 55344 65208 55350
rect 65156 55286 65208 55292
rect 64972 55276 65024 55282
rect 64972 55218 65024 55224
rect 65062 55176 65118 55185
rect 65062 55111 65118 55120
rect 65076 54738 65104 55111
rect 65064 54732 65116 54738
rect 65064 54674 65116 54680
rect 64786 51096 64842 51105
rect 64786 51031 64842 51040
rect 64800 47122 64828 51031
rect 65444 48686 65472 61911
rect 65654 61500 65962 61520
rect 65654 61498 65660 61500
rect 65716 61498 65740 61500
rect 65796 61498 65820 61500
rect 65876 61498 65900 61500
rect 65956 61498 65962 61500
rect 65716 61446 65718 61498
rect 65898 61446 65900 61498
rect 65654 61444 65660 61446
rect 65716 61444 65740 61446
rect 65796 61444 65820 61446
rect 65876 61444 65900 61446
rect 65956 61444 65962 61446
rect 65654 61424 65962 61444
rect 65654 60412 65962 60432
rect 65654 60410 65660 60412
rect 65716 60410 65740 60412
rect 65796 60410 65820 60412
rect 65876 60410 65900 60412
rect 65956 60410 65962 60412
rect 65716 60358 65718 60410
rect 65898 60358 65900 60410
rect 65654 60356 65660 60358
rect 65716 60356 65740 60358
rect 65796 60356 65820 60358
rect 65876 60356 65900 60358
rect 65956 60356 65962 60358
rect 65654 60336 65962 60356
rect 65654 59324 65962 59344
rect 65654 59322 65660 59324
rect 65716 59322 65740 59324
rect 65796 59322 65820 59324
rect 65876 59322 65900 59324
rect 65956 59322 65962 59324
rect 65716 59270 65718 59322
rect 65898 59270 65900 59322
rect 65654 59268 65660 59270
rect 65716 59268 65740 59270
rect 65796 59268 65820 59270
rect 65876 59268 65900 59270
rect 65956 59268 65962 59270
rect 65654 59248 65962 59268
rect 66088 58614 66116 64631
rect 66166 59256 66222 59265
rect 66166 59191 66222 59200
rect 66076 58608 66128 58614
rect 66076 58550 66128 58556
rect 65524 58404 65576 58410
rect 65524 58346 65576 58352
rect 65536 58138 65564 58346
rect 65654 58236 65962 58256
rect 65654 58234 65660 58236
rect 65716 58234 65740 58236
rect 65796 58234 65820 58236
rect 65876 58234 65900 58236
rect 65956 58234 65962 58236
rect 65716 58182 65718 58234
rect 65898 58182 65900 58234
rect 65654 58180 65660 58182
rect 65716 58180 65740 58182
rect 65796 58180 65820 58182
rect 65876 58180 65900 58182
rect 65956 58180 65962 58182
rect 65654 58160 65962 58180
rect 65524 58132 65576 58138
rect 65524 58074 65576 58080
rect 66180 57526 66208 59191
rect 66810 57896 66866 57905
rect 66810 57831 66866 57840
rect 66168 57520 66220 57526
rect 66168 57462 66220 57468
rect 65654 57148 65962 57168
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57072 65962 57092
rect 66166 56536 66222 56545
rect 66166 56471 66222 56480
rect 66180 56234 66208 56471
rect 66168 56228 66220 56234
rect 66168 56170 66220 56176
rect 65654 56060 65962 56080
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55984 65962 56004
rect 66824 55350 66852 57831
rect 66812 55344 66864 55350
rect 66812 55286 66864 55292
rect 65654 54972 65962 54992
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54896 65962 54916
rect 65654 53884 65962 53904
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53808 65962 53828
rect 66074 53816 66130 53825
rect 66074 53751 66130 53760
rect 65654 52796 65962 52816
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52720 65962 52740
rect 65522 52456 65578 52465
rect 65522 52391 65578 52400
rect 65536 51105 65564 52391
rect 65654 51708 65962 51728
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51632 65962 51652
rect 65522 51096 65578 51105
rect 65522 51031 65578 51040
rect 65654 50620 65962 50640
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50544 65962 50564
rect 65654 49532 65962 49552
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49456 65962 49476
rect 65432 48680 65484 48686
rect 65432 48622 65484 48628
rect 65654 48444 65962 48464
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48368 65962 48388
rect 65654 47356 65962 47376
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47280 65962 47300
rect 64788 47116 64840 47122
rect 64788 47058 64840 47064
rect 65654 46268 65962 46288
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46192 65962 46212
rect 65984 45554 66036 45558
rect 66088 45554 66116 53751
rect 66168 47184 66220 47190
rect 66168 47126 66220 47132
rect 66180 47025 66208 47126
rect 66166 47016 66222 47025
rect 66166 46951 66222 46960
rect 65984 45552 66116 45554
rect 66036 45526 66116 45552
rect 65984 45494 66036 45500
rect 65654 45180 65962 45200
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45104 65962 45124
rect 65654 44092 65962 44112
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44016 65962 44036
rect 65654 43004 65962 43024
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42928 65962 42948
rect 66166 42936 66222 42945
rect 66166 42871 66222 42880
rect 66180 42634 66208 42871
rect 66168 42628 66220 42634
rect 66168 42570 66220 42576
rect 65654 41916 65962 41936
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41840 65962 41860
rect 65154 41576 65210 41585
rect 65154 41511 65210 41520
rect 64696 38956 64748 38962
rect 64696 38898 64748 38904
rect 61660 37664 61712 37670
rect 61660 37606 61712 37612
rect 61672 37330 61700 37606
rect 61660 37324 61712 37330
rect 61660 37266 61712 37272
rect 64708 36786 64736 38898
rect 65168 38894 65196 41511
rect 65654 40828 65962 40848
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40752 65962 40772
rect 66166 40216 66222 40225
rect 66166 40151 66222 40160
rect 66180 40118 66208 40151
rect 66168 40112 66220 40118
rect 66168 40054 66220 40060
rect 65654 39740 65962 39760
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39664 65962 39684
rect 65156 38888 65208 38894
rect 65156 38830 65208 38836
rect 65340 38888 65392 38894
rect 67180 38888 67232 38894
rect 65340 38830 65392 38836
rect 67178 38856 67180 38865
rect 67232 38856 67234 38865
rect 65352 38554 65380 38830
rect 67178 38791 67234 38800
rect 65654 38652 65962 38672
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38576 65962 38596
rect 65340 38548 65392 38554
rect 65340 38490 65392 38496
rect 65654 37564 65962 37584
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37488 65962 37508
rect 66166 37496 66222 37505
rect 66166 37431 66222 37440
rect 66180 37330 66208 37431
rect 66168 37324 66220 37330
rect 66168 37266 66220 37272
rect 64696 36780 64748 36786
rect 64696 36722 64748 36728
rect 64880 36576 64932 36582
rect 64880 36518 64932 36524
rect 65524 36576 65576 36582
rect 65524 36518 65576 36524
rect 64892 36310 64920 36518
rect 64880 36304 64932 36310
rect 64880 36246 64932 36252
rect 65536 36242 65564 36518
rect 65654 36476 65962 36496
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36400 65962 36420
rect 65524 36236 65576 36242
rect 65524 36178 65576 36184
rect 67456 36100 67508 36106
rect 67456 36042 67508 36048
rect 61384 35760 61436 35766
rect 61384 35702 61436 35708
rect 61292 35624 61344 35630
rect 61292 35566 61344 35572
rect 59728 30728 59780 30734
rect 59728 30670 59780 30676
rect 60464 30728 60516 30734
rect 60464 30670 60516 30676
rect 59740 29306 59768 30670
rect 60476 30258 60504 30670
rect 60464 30252 60516 30258
rect 60464 30194 60516 30200
rect 59728 29300 59780 29306
rect 59728 29242 59780 29248
rect 60648 28552 60700 28558
rect 60648 28494 60700 28500
rect 60660 28082 60688 28494
rect 60648 28076 60700 28082
rect 60648 28018 60700 28024
rect 60832 28008 60884 28014
rect 60832 27950 60884 27956
rect 60844 27674 60872 27950
rect 60832 27668 60884 27674
rect 60832 27610 60884 27616
rect 61304 27470 61332 35566
rect 65654 35388 65962 35408
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35312 65962 35332
rect 65654 34300 65962 34320
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34224 65962 34244
rect 66076 33584 66128 33590
rect 66076 33526 66128 33532
rect 65654 33212 65962 33232
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33136 65962 33156
rect 65654 32124 65962 32144
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32048 65962 32068
rect 66088 32065 66116 33526
rect 66166 33416 66222 33425
rect 66166 33351 66168 33360
rect 66220 33351 66222 33360
rect 66168 33322 66220 33328
rect 66074 32056 66130 32065
rect 66074 31991 66130 32000
rect 65654 31036 65962 31056
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30960 65962 30980
rect 66166 30696 66222 30705
rect 66166 30631 66168 30640
rect 66220 30631 66222 30640
rect 66168 30602 66220 30608
rect 65654 29948 65962 29968
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29872 65962 29892
rect 61660 29096 61712 29102
rect 61660 29038 61712 29044
rect 61292 27464 61344 27470
rect 61292 27406 61344 27412
rect 58256 26308 58308 26314
rect 58256 26250 58308 26256
rect 58268 26042 58296 26250
rect 58256 26036 58308 26042
rect 58256 25978 58308 25984
rect 58164 25900 58216 25906
rect 58164 25842 58216 25848
rect 57888 22092 57940 22098
rect 57888 22034 57940 22040
rect 57336 3596 57388 3602
rect 57336 3538 57388 3544
rect 57612 3596 57664 3602
rect 57612 3538 57664 3544
rect 57256 3454 57376 3482
rect 57348 800 57376 3454
rect 57900 3398 57928 22034
rect 58176 17678 58204 25842
rect 61672 21554 61700 29038
rect 65654 28860 65962 28880
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28784 65962 28804
rect 64972 28008 65024 28014
rect 64972 27950 65024 27956
rect 66166 27976 66222 27985
rect 64984 25265 65012 27950
rect 66166 27911 66168 27920
rect 66220 27911 66222 27920
rect 66168 27882 66220 27888
rect 65654 27772 65962 27792
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27696 65962 27716
rect 65654 26684 65962 26704
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26608 65962 26628
rect 66166 26616 66222 26625
rect 66166 26551 66222 26560
rect 66180 26382 66208 26551
rect 66168 26376 66220 26382
rect 66168 26318 66220 26324
rect 65654 25596 65962 25616
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25520 65962 25540
rect 64970 25256 65026 25265
rect 64970 25191 65026 25200
rect 65654 24508 65962 24528
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24432 65962 24452
rect 65654 23420 65962 23440
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23344 65962 23364
rect 61752 22432 61804 22438
rect 61752 22374 61804 22380
rect 61764 22098 61792 22374
rect 65654 22332 65962 22352
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22256 65962 22276
rect 61752 22092 61804 22098
rect 61752 22034 61804 22040
rect 61752 21956 61804 21962
rect 61752 21898 61804 21904
rect 66168 21956 66220 21962
rect 66168 21898 66220 21904
rect 61764 21690 61792 21898
rect 66180 21865 66208 21898
rect 66166 21856 66222 21865
rect 66166 21791 66222 21800
rect 61752 21684 61804 21690
rect 61752 21626 61804 21632
rect 61660 21548 61712 21554
rect 61660 21490 61712 21496
rect 61672 20466 61700 21490
rect 65654 21244 65962 21264
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21168 65962 21188
rect 62672 20936 62724 20942
rect 62672 20878 62724 20884
rect 62684 20466 62712 20878
rect 64878 20496 64934 20505
rect 61660 20460 61712 20466
rect 61660 20402 61712 20408
rect 62028 20460 62080 20466
rect 62028 20402 62080 20408
rect 62672 20460 62724 20466
rect 64878 20431 64880 20440
rect 62672 20402 62724 20408
rect 64932 20431 64934 20440
rect 64880 20402 64932 20408
rect 58164 17672 58216 17678
rect 58164 17614 58216 17620
rect 59176 17672 59228 17678
rect 59176 17614 59228 17620
rect 59188 17202 59216 17614
rect 59360 17536 59412 17542
rect 59360 17478 59412 17484
rect 59372 17270 59400 17478
rect 59360 17264 59412 17270
rect 59360 17206 59412 17212
rect 59176 17196 59228 17202
rect 59176 17138 59228 17144
rect 62040 15502 62068 20402
rect 65654 20156 65962 20176
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20080 65962 20100
rect 66168 19304 66220 19310
rect 66168 19246 66220 19252
rect 66180 19145 66208 19246
rect 66166 19136 66222 19145
rect 65654 19068 65962 19088
rect 66166 19071 66222 19080
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 18992 65962 19012
rect 65654 17980 65962 18000
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17904 65962 17924
rect 66168 17876 66220 17882
rect 66168 17818 66220 17824
rect 66180 17785 66208 17818
rect 66166 17776 66222 17785
rect 66166 17711 66222 17720
rect 65524 17128 65576 17134
rect 65524 17070 65576 17076
rect 62028 15496 62080 15502
rect 62028 15438 62080 15444
rect 62856 15496 62908 15502
rect 62856 15438 62908 15444
rect 62868 15026 62896 15438
rect 63224 15360 63276 15366
rect 63224 15302 63276 15308
rect 63236 15094 63264 15302
rect 63224 15088 63276 15094
rect 63224 15030 63276 15036
rect 62856 15020 62908 15026
rect 62856 14962 62908 14968
rect 64788 14952 64840 14958
rect 64788 14894 64840 14900
rect 62120 11688 62172 11694
rect 62120 11630 62172 11636
rect 62132 10674 62160 11630
rect 62120 10668 62172 10674
rect 62120 10610 62172 10616
rect 62764 9988 62816 9994
rect 62764 9930 62816 9936
rect 60648 5160 60700 5166
rect 60648 5102 60700 5108
rect 58624 3596 58676 3602
rect 58624 3538 58676 3544
rect 57888 3392 57940 3398
rect 57888 3334 57940 3340
rect 58636 800 58664 3538
rect 59912 3392 59964 3398
rect 59912 3334 59964 3340
rect 59924 800 59952 3334
rect 60660 2854 60688 5102
rect 62776 4146 62804 9930
rect 64800 4185 64828 14894
rect 64786 4176 64842 4185
rect 62764 4140 62816 4146
rect 64786 4111 64842 4120
rect 62764 4082 62816 4088
rect 65064 3460 65116 3466
rect 65064 3402 65116 3408
rect 60648 2848 60700 2854
rect 60648 2790 60700 2796
rect 63776 2848 63828 2854
rect 63776 2790 63828 2796
rect 63788 800 63816 2790
rect 65076 800 65104 3402
rect 65536 1465 65564 17070
rect 65654 16892 65962 16912
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16816 65962 16836
rect 65654 15804 65962 15824
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15728 65962 15748
rect 65654 14716 65962 14736
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14640 65962 14660
rect 65654 13628 65962 13648
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13552 65962 13572
rect 65654 12540 65962 12560
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12464 65962 12484
rect 65654 11452 65962 11472
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11376 65962 11396
rect 66166 10976 66222 10985
rect 66166 10911 66222 10920
rect 66180 10674 66208 10911
rect 66168 10668 66220 10674
rect 66168 10610 66220 10616
rect 65654 10364 65962 10384
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10288 65962 10308
rect 65654 9276 65962 9296
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9200 65962 9220
rect 66166 8256 66222 8265
rect 65654 8188 65962 8208
rect 66166 8191 66222 8200
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8112 65962 8132
rect 66180 7818 66208 8191
rect 66168 7812 66220 7818
rect 66168 7754 66220 7760
rect 65654 7100 65962 7120
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7024 65962 7044
rect 67468 6914 67496 36042
rect 66824 6886 67496 6914
rect 65654 6012 65962 6032
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5936 65962 5956
rect 65654 4924 65962 4944
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4848 65962 4868
rect 66168 4140 66220 4146
rect 66168 4082 66220 4088
rect 65654 3836 65962 3856
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3760 65962 3780
rect 66180 2825 66208 4082
rect 66166 2816 66222 2825
rect 65654 2748 65962 2768
rect 66166 2751 66222 2760
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2672 65962 2692
rect 65522 1456 65578 1465
rect 65522 1391 65578 1400
rect 66364 870 66576 898
rect 66364 800 66392 870
rect 44652 734 44956 762
rect 45070 0 45182 800
rect 47002 0 47114 800
rect 48290 0 48402 800
rect 49578 0 49690 800
rect 50866 0 50978 800
rect 52154 0 52266 800
rect 53442 0 53554 800
rect 54730 0 54842 800
rect 56018 0 56130 800
rect 57306 0 57418 800
rect 58594 0 58706 800
rect 59882 0 59994 800
rect 61170 0 61282 800
rect 62458 0 62570 800
rect 63746 0 63858 800
rect 65034 0 65146 800
rect 66322 0 66434 800
rect 66548 762 66576 870
rect 66824 762 66852 6886
rect 67640 3664 67692 3670
rect 67640 3606 67692 3612
rect 67652 800 67680 3606
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 68940 800 68968 3470
rect 66548 734 66852 762
rect 67610 0 67722 800
rect 68898 0 69010 800
<< via2 >>
rect 1398 66000 1454 66056
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 3606 68720 3662 68776
rect 3514 67360 3570 67416
rect 3330 64640 3386 64696
rect 3422 61920 3478 61976
rect 3330 59200 3386 59256
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 3698 57840 3754 57896
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3698 46280 3754 46336
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 3422 34040 3478 34096
rect 2962 31320 3018 31376
rect 3422 28600 3478 28656
rect 3146 25880 3202 25936
rect 3422 24520 3478 24576
rect 4066 35400 4122 35456
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 69658 19636 69660
rect 19660 69658 19716 69660
rect 19740 69658 19796 69660
rect 19820 69658 19876 69660
rect 19580 69606 19626 69658
rect 19626 69606 19636 69658
rect 19660 69606 19690 69658
rect 19690 69606 19702 69658
rect 19702 69606 19716 69658
rect 19740 69606 19754 69658
rect 19754 69606 19766 69658
rect 19766 69606 19796 69658
rect 19820 69606 19830 69658
rect 19830 69606 19876 69658
rect 19580 69604 19636 69606
rect 19660 69604 19716 69606
rect 19740 69604 19796 69606
rect 19820 69604 19876 69606
rect 19580 68570 19636 68572
rect 19660 68570 19716 68572
rect 19740 68570 19796 68572
rect 19820 68570 19876 68572
rect 19580 68518 19626 68570
rect 19626 68518 19636 68570
rect 19660 68518 19690 68570
rect 19690 68518 19702 68570
rect 19702 68518 19716 68570
rect 19740 68518 19754 68570
rect 19754 68518 19766 68570
rect 19766 68518 19796 68570
rect 19820 68518 19830 68570
rect 19830 68518 19876 68570
rect 19580 68516 19636 68518
rect 19660 68516 19716 68518
rect 19740 68516 19796 68518
rect 19820 68516 19876 68518
rect 19580 67482 19636 67484
rect 19660 67482 19716 67484
rect 19740 67482 19796 67484
rect 19820 67482 19876 67484
rect 19580 67430 19626 67482
rect 19626 67430 19636 67482
rect 19660 67430 19690 67482
rect 19690 67430 19702 67482
rect 19702 67430 19716 67482
rect 19740 67430 19754 67482
rect 19754 67430 19766 67482
rect 19766 67430 19796 67482
rect 19820 67430 19830 67482
rect 19830 67430 19876 67482
rect 19580 67428 19636 67430
rect 19660 67428 19716 67430
rect 19740 67428 19796 67430
rect 19820 67428 19876 67430
rect 19580 66394 19636 66396
rect 19660 66394 19716 66396
rect 19740 66394 19796 66396
rect 19820 66394 19876 66396
rect 19580 66342 19626 66394
rect 19626 66342 19636 66394
rect 19660 66342 19690 66394
rect 19690 66342 19702 66394
rect 19702 66342 19716 66394
rect 19740 66342 19754 66394
rect 19754 66342 19766 66394
rect 19766 66342 19796 66394
rect 19820 66342 19830 66394
rect 19830 66342 19876 66394
rect 19580 66340 19636 66342
rect 19660 66340 19716 66342
rect 19740 66340 19796 66342
rect 19820 66340 19876 66342
rect 19580 65306 19636 65308
rect 19660 65306 19716 65308
rect 19740 65306 19796 65308
rect 19820 65306 19876 65308
rect 19580 65254 19626 65306
rect 19626 65254 19636 65306
rect 19660 65254 19690 65306
rect 19690 65254 19702 65306
rect 19702 65254 19716 65306
rect 19740 65254 19754 65306
rect 19754 65254 19766 65306
rect 19766 65254 19796 65306
rect 19820 65254 19830 65306
rect 19830 65254 19876 65306
rect 19580 65252 19636 65254
rect 19660 65252 19716 65254
rect 19740 65252 19796 65254
rect 19820 65252 19876 65254
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4066 21836 4068 21856
rect 4068 21836 4120 21856
rect 4120 21836 4122 21856
rect 4066 21800 4122 21836
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4066 20440 4122 20496
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4066 16396 4068 16416
rect 4068 16396 4120 16416
rect 4120 16396 4122 16416
rect 4066 16360 4122 16396
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 3974 15000 4030 15056
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4066 13640 4122 13696
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3422 10956 3424 10976
rect 3424 10956 3476 10976
rect 3476 10956 3478 10976
rect 3422 10920 3478 10956
rect 3422 9596 3424 9616
rect 3424 9596 3476 9616
rect 3476 9596 3478 9616
rect 3422 9560 3478 9596
rect 3422 8236 3424 8256
rect 3424 8236 3476 8256
rect 3476 8236 3478 8256
rect 3422 8200 3478 8236
rect 3422 6840 3478 6896
rect 3422 5480 3478 5536
rect 3146 4120 3202 4176
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3514 2760 3570 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 64218 19636 64220
rect 19660 64218 19716 64220
rect 19740 64218 19796 64220
rect 19820 64218 19876 64220
rect 19580 64166 19626 64218
rect 19626 64166 19636 64218
rect 19660 64166 19690 64218
rect 19690 64166 19702 64218
rect 19702 64166 19716 64218
rect 19740 64166 19754 64218
rect 19754 64166 19766 64218
rect 19766 64166 19796 64218
rect 19820 64166 19830 64218
rect 19830 64166 19876 64218
rect 19580 64164 19636 64166
rect 19660 64164 19716 64166
rect 19740 64164 19796 64166
rect 19820 64164 19876 64166
rect 19580 63130 19636 63132
rect 19660 63130 19716 63132
rect 19740 63130 19796 63132
rect 19820 63130 19876 63132
rect 19580 63078 19626 63130
rect 19626 63078 19636 63130
rect 19660 63078 19690 63130
rect 19690 63078 19702 63130
rect 19702 63078 19716 63130
rect 19740 63078 19754 63130
rect 19754 63078 19766 63130
rect 19766 63078 19796 63130
rect 19820 63078 19830 63130
rect 19830 63078 19876 63130
rect 19580 63076 19636 63078
rect 19660 63076 19716 63078
rect 19740 63076 19796 63078
rect 19820 63076 19876 63078
rect 19580 62042 19636 62044
rect 19660 62042 19716 62044
rect 19740 62042 19796 62044
rect 19820 62042 19876 62044
rect 19580 61990 19626 62042
rect 19626 61990 19636 62042
rect 19660 61990 19690 62042
rect 19690 61990 19702 62042
rect 19702 61990 19716 62042
rect 19740 61990 19754 62042
rect 19754 61990 19766 62042
rect 19766 61990 19796 62042
rect 19820 61990 19830 62042
rect 19830 61990 19876 62042
rect 19580 61988 19636 61990
rect 19660 61988 19716 61990
rect 19740 61988 19796 61990
rect 19820 61988 19876 61990
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 34940 69114 34996 69116
rect 35020 69114 35076 69116
rect 35100 69114 35156 69116
rect 35180 69114 35236 69116
rect 34940 69062 34986 69114
rect 34986 69062 34996 69114
rect 35020 69062 35050 69114
rect 35050 69062 35062 69114
rect 35062 69062 35076 69114
rect 35100 69062 35114 69114
rect 35114 69062 35126 69114
rect 35126 69062 35156 69114
rect 35180 69062 35190 69114
rect 35190 69062 35236 69114
rect 34940 69060 34996 69062
rect 35020 69060 35076 69062
rect 35100 69060 35156 69062
rect 35180 69060 35236 69062
rect 34940 68026 34996 68028
rect 35020 68026 35076 68028
rect 35100 68026 35156 68028
rect 35180 68026 35236 68028
rect 34940 67974 34986 68026
rect 34986 67974 34996 68026
rect 35020 67974 35050 68026
rect 35050 67974 35062 68026
rect 35062 67974 35076 68026
rect 35100 67974 35114 68026
rect 35114 67974 35126 68026
rect 35126 67974 35156 68026
rect 35180 67974 35190 68026
rect 35190 67974 35236 68026
rect 34940 67972 34996 67974
rect 35020 67972 35076 67974
rect 35100 67972 35156 67974
rect 35180 67972 35236 67974
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 34940 64762 34996 64764
rect 35020 64762 35076 64764
rect 35100 64762 35156 64764
rect 35180 64762 35236 64764
rect 34940 64710 34986 64762
rect 34986 64710 34996 64762
rect 35020 64710 35050 64762
rect 35050 64710 35062 64762
rect 35062 64710 35076 64762
rect 35100 64710 35114 64762
rect 35114 64710 35126 64762
rect 35126 64710 35156 64762
rect 35180 64710 35190 64762
rect 35190 64710 35236 64762
rect 34940 64708 34996 64710
rect 35020 64708 35076 64710
rect 35100 64708 35156 64710
rect 35180 64708 35236 64710
rect 34940 63674 34996 63676
rect 35020 63674 35076 63676
rect 35100 63674 35156 63676
rect 35180 63674 35236 63676
rect 34940 63622 34986 63674
rect 34986 63622 34996 63674
rect 35020 63622 35050 63674
rect 35050 63622 35062 63674
rect 35062 63622 35076 63674
rect 35100 63622 35114 63674
rect 35114 63622 35126 63674
rect 35126 63622 35156 63674
rect 35180 63622 35190 63674
rect 35190 63622 35236 63674
rect 34940 63620 34996 63622
rect 35020 63620 35076 63622
rect 35100 63620 35156 63622
rect 35180 63620 35236 63622
rect 34940 62586 34996 62588
rect 35020 62586 35076 62588
rect 35100 62586 35156 62588
rect 35180 62586 35236 62588
rect 34940 62534 34986 62586
rect 34986 62534 34996 62586
rect 35020 62534 35050 62586
rect 35050 62534 35062 62586
rect 35062 62534 35076 62586
rect 35100 62534 35114 62586
rect 35114 62534 35126 62586
rect 35126 62534 35156 62586
rect 35180 62534 35190 62586
rect 35190 62534 35236 62586
rect 34940 62532 34996 62534
rect 35020 62532 35076 62534
rect 35100 62532 35156 62534
rect 35180 62532 35236 62534
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 69658 50356 69660
rect 50380 69658 50436 69660
rect 50460 69658 50516 69660
rect 50540 69658 50596 69660
rect 50300 69606 50346 69658
rect 50346 69606 50356 69658
rect 50380 69606 50410 69658
rect 50410 69606 50422 69658
rect 50422 69606 50436 69658
rect 50460 69606 50474 69658
rect 50474 69606 50486 69658
rect 50486 69606 50516 69658
rect 50540 69606 50550 69658
rect 50550 69606 50596 69658
rect 50300 69604 50356 69606
rect 50380 69604 50436 69606
rect 50460 69604 50516 69606
rect 50540 69604 50596 69606
rect 50300 68570 50356 68572
rect 50380 68570 50436 68572
rect 50460 68570 50516 68572
rect 50540 68570 50596 68572
rect 50300 68518 50346 68570
rect 50346 68518 50356 68570
rect 50380 68518 50410 68570
rect 50410 68518 50422 68570
rect 50422 68518 50436 68570
rect 50460 68518 50474 68570
rect 50474 68518 50486 68570
rect 50486 68518 50516 68570
rect 50540 68518 50550 68570
rect 50550 68518 50596 68570
rect 50300 68516 50356 68518
rect 50380 68516 50436 68518
rect 50460 68516 50516 68518
rect 50540 68516 50596 68518
rect 50300 67482 50356 67484
rect 50380 67482 50436 67484
rect 50460 67482 50516 67484
rect 50540 67482 50596 67484
rect 50300 67430 50346 67482
rect 50346 67430 50356 67482
rect 50380 67430 50410 67482
rect 50410 67430 50422 67482
rect 50422 67430 50436 67482
rect 50460 67430 50474 67482
rect 50474 67430 50486 67482
rect 50486 67430 50516 67482
rect 50540 67430 50550 67482
rect 50550 67430 50596 67482
rect 50300 67428 50356 67430
rect 50380 67428 50436 67430
rect 50460 67428 50516 67430
rect 50540 67428 50596 67430
rect 50300 66394 50356 66396
rect 50380 66394 50436 66396
rect 50460 66394 50516 66396
rect 50540 66394 50596 66396
rect 50300 66342 50346 66394
rect 50346 66342 50356 66394
rect 50380 66342 50410 66394
rect 50410 66342 50422 66394
rect 50422 66342 50436 66394
rect 50460 66342 50474 66394
rect 50474 66342 50486 66394
rect 50486 66342 50516 66394
rect 50540 66342 50550 66394
rect 50550 66342 50596 66394
rect 50300 66340 50356 66342
rect 50380 66340 50436 66342
rect 50460 66340 50516 66342
rect 50540 66340 50596 66342
rect 50300 65306 50356 65308
rect 50380 65306 50436 65308
rect 50460 65306 50516 65308
rect 50540 65306 50596 65308
rect 50300 65254 50346 65306
rect 50346 65254 50356 65306
rect 50380 65254 50410 65306
rect 50410 65254 50422 65306
rect 50422 65254 50436 65306
rect 50460 65254 50474 65306
rect 50474 65254 50486 65306
rect 50486 65254 50516 65306
rect 50540 65254 50550 65306
rect 50550 65254 50596 65306
rect 50300 65252 50356 65254
rect 50380 65252 50436 65254
rect 50460 65252 50516 65254
rect 50540 65252 50596 65254
rect 50300 64218 50356 64220
rect 50380 64218 50436 64220
rect 50460 64218 50516 64220
rect 50540 64218 50596 64220
rect 50300 64166 50346 64218
rect 50346 64166 50356 64218
rect 50380 64166 50410 64218
rect 50410 64166 50422 64218
rect 50422 64166 50436 64218
rect 50460 64166 50474 64218
rect 50474 64166 50486 64218
rect 50486 64166 50516 64218
rect 50540 64166 50550 64218
rect 50550 64166 50596 64218
rect 50300 64164 50356 64166
rect 50380 64164 50436 64166
rect 50460 64164 50516 64166
rect 50540 64164 50596 64166
rect 50300 63130 50356 63132
rect 50380 63130 50436 63132
rect 50460 63130 50516 63132
rect 50540 63130 50596 63132
rect 50300 63078 50346 63130
rect 50346 63078 50356 63130
rect 50380 63078 50410 63130
rect 50410 63078 50422 63130
rect 50422 63078 50436 63130
rect 50460 63078 50474 63130
rect 50474 63078 50486 63130
rect 50486 63078 50516 63130
rect 50540 63078 50550 63130
rect 50550 63078 50596 63130
rect 50300 63076 50356 63078
rect 50380 63076 50436 63078
rect 50460 63076 50516 63078
rect 50540 63076 50596 63078
rect 50300 62042 50356 62044
rect 50380 62042 50436 62044
rect 50460 62042 50516 62044
rect 50540 62042 50596 62044
rect 50300 61990 50346 62042
rect 50346 61990 50356 62042
rect 50380 61990 50410 62042
rect 50410 61990 50422 62042
rect 50422 61990 50436 62042
rect 50460 61990 50474 62042
rect 50474 61990 50486 62042
rect 50486 61990 50516 62042
rect 50540 61990 50550 62042
rect 50550 61990 50596 62042
rect 50300 61988 50356 61990
rect 50380 61988 50436 61990
rect 50460 61988 50516 61990
rect 50540 61988 50596 61990
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 66074 70080 66130 70136
rect 65660 69114 65716 69116
rect 65740 69114 65796 69116
rect 65820 69114 65876 69116
rect 65900 69114 65956 69116
rect 65660 69062 65706 69114
rect 65706 69062 65716 69114
rect 65740 69062 65770 69114
rect 65770 69062 65782 69114
rect 65782 69062 65796 69114
rect 65820 69062 65834 69114
rect 65834 69062 65846 69114
rect 65846 69062 65876 69114
rect 65900 69062 65910 69114
rect 65910 69062 65956 69114
rect 65660 69060 65716 69062
rect 65740 69060 65796 69062
rect 65820 69060 65876 69062
rect 65900 69060 65956 69062
rect 65660 68026 65716 68028
rect 65740 68026 65796 68028
rect 65820 68026 65876 68028
rect 65900 68026 65956 68028
rect 65660 67974 65706 68026
rect 65706 67974 65716 68026
rect 65740 67974 65770 68026
rect 65770 67974 65782 68026
rect 65782 67974 65796 68026
rect 65820 67974 65834 68026
rect 65834 67974 65846 68026
rect 65846 67974 65876 68026
rect 65900 67974 65910 68026
rect 65910 67974 65956 68026
rect 65660 67972 65716 67974
rect 65740 67972 65796 67974
rect 65820 67972 65876 67974
rect 65900 67972 65956 67974
rect 65338 67360 65394 67416
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 64878 66000 64934 66056
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 65660 64762 65716 64764
rect 65740 64762 65796 64764
rect 65820 64762 65876 64764
rect 65900 64762 65956 64764
rect 65660 64710 65706 64762
rect 65706 64710 65716 64762
rect 65740 64710 65770 64762
rect 65770 64710 65782 64762
rect 65782 64710 65796 64762
rect 65820 64710 65834 64762
rect 65834 64710 65846 64762
rect 65846 64710 65876 64762
rect 65900 64710 65910 64762
rect 65910 64710 65956 64762
rect 65660 64708 65716 64710
rect 65740 64708 65796 64710
rect 65820 64708 65876 64710
rect 65900 64708 65956 64710
rect 66074 64640 66130 64696
rect 65660 63674 65716 63676
rect 65740 63674 65796 63676
rect 65820 63674 65876 63676
rect 65900 63674 65956 63676
rect 65660 63622 65706 63674
rect 65706 63622 65716 63674
rect 65740 63622 65770 63674
rect 65770 63622 65782 63674
rect 65782 63622 65796 63674
rect 65820 63622 65834 63674
rect 65834 63622 65846 63674
rect 65846 63622 65876 63674
rect 65900 63622 65910 63674
rect 65910 63622 65956 63674
rect 65660 63620 65716 63622
rect 65740 63620 65796 63622
rect 65820 63620 65876 63622
rect 65900 63620 65956 63622
rect 65660 62586 65716 62588
rect 65740 62586 65796 62588
rect 65820 62586 65876 62588
rect 65900 62586 65956 62588
rect 65660 62534 65706 62586
rect 65706 62534 65716 62586
rect 65740 62534 65770 62586
rect 65770 62534 65782 62586
rect 65782 62534 65796 62586
rect 65820 62534 65834 62586
rect 65834 62534 65846 62586
rect 65846 62534 65876 62586
rect 65900 62534 65910 62586
rect 65910 62534 65956 62586
rect 65660 62532 65716 62534
rect 65740 62532 65796 62534
rect 65820 62532 65876 62534
rect 65900 62532 65956 62534
rect 65430 61920 65486 61976
rect 65062 55120 65118 55176
rect 64786 51040 64842 51096
rect 65660 61498 65716 61500
rect 65740 61498 65796 61500
rect 65820 61498 65876 61500
rect 65900 61498 65956 61500
rect 65660 61446 65706 61498
rect 65706 61446 65716 61498
rect 65740 61446 65770 61498
rect 65770 61446 65782 61498
rect 65782 61446 65796 61498
rect 65820 61446 65834 61498
rect 65834 61446 65846 61498
rect 65846 61446 65876 61498
rect 65900 61446 65910 61498
rect 65910 61446 65956 61498
rect 65660 61444 65716 61446
rect 65740 61444 65796 61446
rect 65820 61444 65876 61446
rect 65900 61444 65956 61446
rect 65660 60410 65716 60412
rect 65740 60410 65796 60412
rect 65820 60410 65876 60412
rect 65900 60410 65956 60412
rect 65660 60358 65706 60410
rect 65706 60358 65716 60410
rect 65740 60358 65770 60410
rect 65770 60358 65782 60410
rect 65782 60358 65796 60410
rect 65820 60358 65834 60410
rect 65834 60358 65846 60410
rect 65846 60358 65876 60410
rect 65900 60358 65910 60410
rect 65910 60358 65956 60410
rect 65660 60356 65716 60358
rect 65740 60356 65796 60358
rect 65820 60356 65876 60358
rect 65900 60356 65956 60358
rect 65660 59322 65716 59324
rect 65740 59322 65796 59324
rect 65820 59322 65876 59324
rect 65900 59322 65956 59324
rect 65660 59270 65706 59322
rect 65706 59270 65716 59322
rect 65740 59270 65770 59322
rect 65770 59270 65782 59322
rect 65782 59270 65796 59322
rect 65820 59270 65834 59322
rect 65834 59270 65846 59322
rect 65846 59270 65876 59322
rect 65900 59270 65910 59322
rect 65910 59270 65956 59322
rect 65660 59268 65716 59270
rect 65740 59268 65796 59270
rect 65820 59268 65876 59270
rect 65900 59268 65956 59270
rect 66166 59200 66222 59256
rect 65660 58234 65716 58236
rect 65740 58234 65796 58236
rect 65820 58234 65876 58236
rect 65900 58234 65956 58236
rect 65660 58182 65706 58234
rect 65706 58182 65716 58234
rect 65740 58182 65770 58234
rect 65770 58182 65782 58234
rect 65782 58182 65796 58234
rect 65820 58182 65834 58234
rect 65834 58182 65846 58234
rect 65846 58182 65876 58234
rect 65900 58182 65910 58234
rect 65910 58182 65956 58234
rect 65660 58180 65716 58182
rect 65740 58180 65796 58182
rect 65820 58180 65876 58182
rect 65900 58180 65956 58182
rect 66810 57840 66866 57896
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 66166 56480 66222 56536
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 66074 53760 66130 53816
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 65522 52400 65578 52456
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 65522 51040 65578 51096
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 66166 46960 66222 47016
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 66166 42880 66222 42936
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 65154 41520 65210 41576
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 66166 40160 66222 40216
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 67178 38836 67180 38856
rect 67180 38836 67232 38856
rect 67232 38836 67234 38856
rect 67178 38800 67234 38836
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 66166 37440 66222 37496
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 66166 33380 66222 33416
rect 66166 33360 66168 33380
rect 66168 33360 66220 33380
rect 66220 33360 66222 33380
rect 66074 32000 66130 32056
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 66166 30660 66222 30696
rect 66166 30640 66168 30660
rect 66168 30640 66220 30660
rect 66220 30640 66222 30660
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 66166 27940 66222 27976
rect 66166 27920 66168 27940
rect 66168 27920 66220 27940
rect 66220 27920 66222 27940
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 66166 26560 66222 26616
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 64970 25200 65026 25256
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 66166 21800 66222 21856
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 64878 20460 64934 20496
rect 64878 20440 64880 20460
rect 64880 20440 64932 20460
rect 64932 20440 64934 20460
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 66166 19080 66222 19136
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 66166 17720 66222 17776
rect 64786 4120 64842 4176
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 66166 10920 66222 10976
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 66166 8200 66222 8256
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 66166 2760 66222 2816
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 65522 1400 65578 1456
<< metal3 >>
rect 0 71348 800 71588
rect 0 69988 800 70228
rect 66069 70138 66135 70141
rect 69200 70138 70000 70228
rect 66069 70136 70000 70138
rect 66069 70080 66074 70136
rect 66130 70080 70000 70136
rect 66069 70078 70000 70080
rect 66069 70075 66135 70078
rect 69200 69988 70000 70078
rect 19568 69664 19888 69665
rect 19568 69600 19576 69664
rect 19640 69600 19656 69664
rect 19720 69600 19736 69664
rect 19800 69600 19816 69664
rect 19880 69600 19888 69664
rect 19568 69599 19888 69600
rect 50288 69664 50608 69665
rect 50288 69600 50296 69664
rect 50360 69600 50376 69664
rect 50440 69600 50456 69664
rect 50520 69600 50536 69664
rect 50600 69600 50608 69664
rect 50288 69599 50608 69600
rect 4208 69120 4528 69121
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 69055 4528 69056
rect 34928 69120 35248 69121
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 69055 35248 69056
rect 65648 69120 65968 69121
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 69055 65968 69056
rect 0 68778 800 68868
rect 3601 68778 3667 68781
rect 0 68776 3667 68778
rect 0 68720 3606 68776
rect 3662 68720 3667 68776
rect 0 68718 3667 68720
rect 0 68628 800 68718
rect 3601 68715 3667 68718
rect 69200 68628 70000 68868
rect 19568 68576 19888 68577
rect 19568 68512 19576 68576
rect 19640 68512 19656 68576
rect 19720 68512 19736 68576
rect 19800 68512 19816 68576
rect 19880 68512 19888 68576
rect 19568 68511 19888 68512
rect 50288 68576 50608 68577
rect 50288 68512 50296 68576
rect 50360 68512 50376 68576
rect 50440 68512 50456 68576
rect 50520 68512 50536 68576
rect 50600 68512 50608 68576
rect 50288 68511 50608 68512
rect 4208 68032 4528 68033
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 67967 4528 67968
rect 34928 68032 35248 68033
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 67967 35248 67968
rect 65648 68032 65968 68033
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 67967 65968 67968
rect 0 67418 800 67508
rect 19568 67488 19888 67489
rect 19568 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19888 67488
rect 19568 67423 19888 67424
rect 50288 67488 50608 67489
rect 50288 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50608 67488
rect 50288 67423 50608 67424
rect 3509 67418 3575 67421
rect 0 67416 3575 67418
rect 0 67360 3514 67416
rect 3570 67360 3575 67416
rect 0 67358 3575 67360
rect 0 67268 800 67358
rect 3509 67355 3575 67358
rect 65333 67418 65399 67421
rect 69200 67418 70000 67508
rect 65333 67416 70000 67418
rect 65333 67360 65338 67416
rect 65394 67360 70000 67416
rect 65333 67358 70000 67360
rect 65333 67355 65399 67358
rect 69200 67268 70000 67358
rect 4208 66944 4528 66945
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 66879 4528 66880
rect 34928 66944 35248 66945
rect 34928 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35248 66944
rect 34928 66879 35248 66880
rect 65648 66944 65968 66945
rect 65648 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65968 66944
rect 65648 66879 65968 66880
rect 19568 66400 19888 66401
rect 19568 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19888 66400
rect 19568 66335 19888 66336
rect 50288 66400 50608 66401
rect 50288 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50608 66400
rect 50288 66335 50608 66336
rect 0 66058 800 66148
rect 1393 66058 1459 66061
rect 0 66056 1459 66058
rect 0 66000 1398 66056
rect 1454 66000 1459 66056
rect 0 65998 1459 66000
rect 0 65908 800 65998
rect 1393 65995 1459 65998
rect 64873 66058 64939 66061
rect 69200 66058 70000 66148
rect 64873 66056 70000 66058
rect 64873 66000 64878 66056
rect 64934 66000 70000 66056
rect 64873 65998 70000 66000
rect 64873 65995 64939 65998
rect 69200 65908 70000 65998
rect 4208 65856 4528 65857
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 65791 4528 65792
rect 34928 65856 35248 65857
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 65791 35248 65792
rect 65648 65856 65968 65857
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 65791 65968 65792
rect 19568 65312 19888 65313
rect 19568 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19888 65312
rect 19568 65247 19888 65248
rect 50288 65312 50608 65313
rect 50288 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50608 65312
rect 50288 65247 50608 65248
rect 0 64698 800 64788
rect 4208 64768 4528 64769
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 64703 4528 64704
rect 34928 64768 35248 64769
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 64703 35248 64704
rect 65648 64768 65968 64769
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 64703 65968 64704
rect 3325 64698 3391 64701
rect 0 64696 3391 64698
rect 0 64640 3330 64696
rect 3386 64640 3391 64696
rect 0 64638 3391 64640
rect 0 64548 800 64638
rect 3325 64635 3391 64638
rect 66069 64698 66135 64701
rect 69200 64698 70000 64788
rect 66069 64696 70000 64698
rect 66069 64640 66074 64696
rect 66130 64640 70000 64696
rect 66069 64638 70000 64640
rect 66069 64635 66135 64638
rect 69200 64548 70000 64638
rect 19568 64224 19888 64225
rect 19568 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19888 64224
rect 19568 64159 19888 64160
rect 50288 64224 50608 64225
rect 50288 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50608 64224
rect 50288 64159 50608 64160
rect 4208 63680 4528 63681
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 63615 4528 63616
rect 34928 63680 35248 63681
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 63615 35248 63616
rect 65648 63680 65968 63681
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 63615 65968 63616
rect 0 63188 800 63428
rect 69200 63188 70000 63428
rect 19568 63136 19888 63137
rect 19568 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19888 63136
rect 19568 63071 19888 63072
rect 50288 63136 50608 63137
rect 50288 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50608 63136
rect 50288 63071 50608 63072
rect 4208 62592 4528 62593
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 62527 4528 62528
rect 34928 62592 35248 62593
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 62527 35248 62528
rect 65648 62592 65968 62593
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 62527 65968 62528
rect 0 61978 800 62068
rect 19568 62048 19888 62049
rect 19568 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19888 62048
rect 19568 61983 19888 61984
rect 50288 62048 50608 62049
rect 50288 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50608 62048
rect 50288 61983 50608 61984
rect 3417 61978 3483 61981
rect 0 61976 3483 61978
rect 0 61920 3422 61976
rect 3478 61920 3483 61976
rect 0 61918 3483 61920
rect 0 61828 800 61918
rect 3417 61915 3483 61918
rect 65425 61978 65491 61981
rect 69200 61978 70000 62068
rect 65425 61976 70000 61978
rect 65425 61920 65430 61976
rect 65486 61920 70000 61976
rect 65425 61918 70000 61920
rect 65425 61915 65491 61918
rect 69200 61828 70000 61918
rect 4208 61504 4528 61505
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 61439 4528 61440
rect 34928 61504 35248 61505
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 61439 35248 61440
rect 65648 61504 65968 61505
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 61439 65968 61440
rect 19568 60960 19888 60961
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 60895 19888 60896
rect 50288 60960 50608 60961
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 60895 50608 60896
rect 0 60468 800 60708
rect 69200 60468 70000 60708
rect 4208 60416 4528 60417
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 60351 4528 60352
rect 34928 60416 35248 60417
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 60351 35248 60352
rect 65648 60416 65968 60417
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 60351 65968 60352
rect 19568 59872 19888 59873
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 59807 19888 59808
rect 50288 59872 50608 59873
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 59807 50608 59808
rect 0 59258 800 59348
rect 4208 59328 4528 59329
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 59263 4528 59264
rect 34928 59328 35248 59329
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 59263 35248 59264
rect 65648 59328 65968 59329
rect 65648 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65968 59328
rect 65648 59263 65968 59264
rect 3325 59258 3391 59261
rect 0 59256 3391 59258
rect 0 59200 3330 59256
rect 3386 59200 3391 59256
rect 0 59198 3391 59200
rect 0 59108 800 59198
rect 3325 59195 3391 59198
rect 66161 59258 66227 59261
rect 69200 59258 70000 59348
rect 66161 59256 70000 59258
rect 66161 59200 66166 59256
rect 66222 59200 70000 59256
rect 66161 59198 70000 59200
rect 66161 59195 66227 59198
rect 69200 59108 70000 59198
rect 19568 58784 19888 58785
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 58719 19888 58720
rect 50288 58784 50608 58785
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 58719 50608 58720
rect 4208 58240 4528 58241
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 58175 4528 58176
rect 34928 58240 35248 58241
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 58175 35248 58176
rect 65648 58240 65968 58241
rect 65648 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65968 58240
rect 65648 58175 65968 58176
rect 0 57898 800 57988
rect 3693 57898 3759 57901
rect 0 57896 3759 57898
rect 0 57840 3698 57896
rect 3754 57840 3759 57896
rect 0 57838 3759 57840
rect 0 57748 800 57838
rect 3693 57835 3759 57838
rect 66805 57898 66871 57901
rect 69200 57898 70000 57988
rect 66805 57896 70000 57898
rect 66805 57840 66810 57896
rect 66866 57840 70000 57896
rect 66805 57838 70000 57840
rect 66805 57835 66871 57838
rect 69200 57748 70000 57838
rect 19568 57696 19888 57697
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 57631 19888 57632
rect 50288 57696 50608 57697
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 57631 50608 57632
rect 4208 57152 4528 57153
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 57087 4528 57088
rect 34928 57152 35248 57153
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 57087 35248 57088
rect 65648 57152 65968 57153
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 57087 65968 57088
rect 0 56388 800 56628
rect 19568 56608 19888 56609
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 56543 19888 56544
rect 50288 56608 50608 56609
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 56543 50608 56544
rect 66161 56538 66227 56541
rect 69200 56538 70000 56628
rect 66161 56536 70000 56538
rect 66161 56480 66166 56536
rect 66222 56480 70000 56536
rect 66161 56478 70000 56480
rect 66161 56475 66227 56478
rect 69200 56388 70000 56478
rect 4208 56064 4528 56065
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 55999 4528 56000
rect 34928 56064 35248 56065
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 55999 35248 56000
rect 65648 56064 65968 56065
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 55999 65968 56000
rect 19568 55520 19888 55521
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 55455 19888 55456
rect 50288 55520 50608 55521
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 55455 50608 55456
rect 0 55028 800 55268
rect 65057 55178 65123 55181
rect 69200 55178 70000 55268
rect 65057 55176 70000 55178
rect 65057 55120 65062 55176
rect 65118 55120 70000 55176
rect 65057 55118 70000 55120
rect 65057 55115 65123 55118
rect 69200 55028 70000 55118
rect 4208 54976 4528 54977
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 54911 4528 54912
rect 34928 54976 35248 54977
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 54911 35248 54912
rect 65648 54976 65968 54977
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 54911 65968 54912
rect 19568 54432 19888 54433
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 54367 19888 54368
rect 50288 54432 50608 54433
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 54367 50608 54368
rect 0 53668 800 53908
rect 4208 53888 4528 53889
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 53823 4528 53824
rect 34928 53888 35248 53889
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 53823 35248 53824
rect 65648 53888 65968 53889
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 53823 65968 53824
rect 66069 53818 66135 53821
rect 69200 53818 70000 53908
rect 66069 53816 70000 53818
rect 66069 53760 66074 53816
rect 66130 53760 70000 53816
rect 66069 53758 70000 53760
rect 66069 53755 66135 53758
rect 69200 53668 70000 53758
rect 19568 53344 19888 53345
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 53279 19888 53280
rect 50288 53344 50608 53345
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 53279 50608 53280
rect 4208 52800 4528 52801
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 52735 4528 52736
rect 34928 52800 35248 52801
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 52735 35248 52736
rect 65648 52800 65968 52801
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 52735 65968 52736
rect 0 52308 800 52548
rect 65517 52458 65583 52461
rect 69200 52458 70000 52548
rect 65517 52456 70000 52458
rect 65517 52400 65522 52456
rect 65578 52400 70000 52456
rect 65517 52398 70000 52400
rect 65517 52395 65583 52398
rect 69200 52308 70000 52398
rect 19568 52256 19888 52257
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 52191 19888 52192
rect 50288 52256 50608 52257
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 52191 50608 52192
rect 4208 51712 4528 51713
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 51647 4528 51648
rect 34928 51712 35248 51713
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 51647 35248 51648
rect 65648 51712 65968 51713
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 51647 65968 51648
rect 0 50948 800 51188
rect 19568 51168 19888 51169
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 51103 19888 51104
rect 50288 51168 50608 51169
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 51103 50608 51104
rect 64781 51098 64847 51101
rect 65517 51098 65583 51101
rect 64781 51096 65583 51098
rect 64781 51040 64786 51096
rect 64842 51040 65522 51096
rect 65578 51040 65583 51096
rect 64781 51038 65583 51040
rect 64781 51035 64847 51038
rect 65517 51035 65583 51038
rect 69200 50948 70000 51188
rect 4208 50624 4528 50625
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 50559 4528 50560
rect 34928 50624 35248 50625
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 50559 35248 50560
rect 65648 50624 65968 50625
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 50559 65968 50560
rect 19568 50080 19888 50081
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 50015 19888 50016
rect 50288 50080 50608 50081
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 50015 50608 50016
rect 0 49588 800 49828
rect 69200 49588 70000 49828
rect 4208 49536 4528 49537
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 49471 4528 49472
rect 34928 49536 35248 49537
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 49471 35248 49472
rect 65648 49536 65968 49537
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 49471 65968 49472
rect 19568 48992 19888 48993
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 48927 19888 48928
rect 50288 48992 50608 48993
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 48927 50608 48928
rect 4208 48448 4528 48449
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 48383 4528 48384
rect 34928 48448 35248 48449
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 48383 35248 48384
rect 65648 48448 65968 48449
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 48383 65968 48384
rect 69200 48228 70000 48468
rect 19568 47904 19888 47905
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 47839 19888 47840
rect 50288 47904 50608 47905
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 47839 50608 47840
rect 0 47548 800 47788
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 65648 47360 65968 47361
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 47295 65968 47296
rect 66161 47018 66227 47021
rect 69200 47018 70000 47108
rect 66161 47016 70000 47018
rect 66161 46960 66166 47016
rect 66222 46960 70000 47016
rect 66161 46958 70000 46960
rect 66161 46955 66227 46958
rect 69200 46868 70000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 50288 46816 50608 46817
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 46751 50608 46752
rect 0 46338 800 46428
rect 3693 46338 3759 46341
rect 0 46336 3759 46338
rect 0 46280 3698 46336
rect 3754 46280 3759 46336
rect 0 46278 3759 46280
rect 0 46188 800 46278
rect 3693 46275 3759 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 65648 46272 65968 46273
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 46207 65968 46208
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 50288 45728 50608 45729
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 45663 50608 45664
rect 69200 45508 70000 45748
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 65648 45184 65968 45185
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 45119 65968 45120
rect 0 44828 800 45068
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 50288 44640 50608 44641
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 44575 50608 44576
rect 69200 44148 70000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 65648 44096 65968 44097
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 44031 65968 44032
rect 0 43468 800 43708
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 50288 43552 50608 43553
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 43487 50608 43488
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 65648 43008 65968 43009
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 42943 65968 42944
rect 66161 42938 66227 42941
rect 69200 42938 70000 43028
rect 66161 42936 70000 42938
rect 66161 42880 66166 42936
rect 66222 42880 70000 42936
rect 66161 42878 70000 42880
rect 66161 42875 66227 42878
rect 69200 42788 70000 42878
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 50288 42464 50608 42465
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 42399 50608 42400
rect 0 42108 800 42348
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 65648 41920 65968 41921
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 41855 65968 41856
rect 65149 41578 65215 41581
rect 69200 41578 70000 41668
rect 65149 41576 70000 41578
rect 65149 41520 65154 41576
rect 65210 41520 70000 41576
rect 65149 41518 70000 41520
rect 65149 41515 65215 41518
rect 69200 41428 70000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 50288 41376 50608 41377
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 41311 50608 41312
rect 0 40748 800 40988
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 65648 40832 65968 40833
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 40767 65968 40768
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 50288 40288 50608 40289
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 40223 50608 40224
rect 66161 40218 66227 40221
rect 69200 40218 70000 40308
rect 66161 40216 70000 40218
rect 66161 40160 66166 40216
rect 66222 40160 70000 40216
rect 66161 40158 70000 40160
rect 66161 40155 66227 40158
rect 69200 40068 70000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 65648 39744 65968 39745
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 39679 65968 39680
rect 0 39388 800 39628
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 50288 39200 50608 39201
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 39135 50608 39136
rect 67173 38858 67239 38861
rect 69200 38858 70000 38948
rect 67173 38856 70000 38858
rect 67173 38800 67178 38856
rect 67234 38800 70000 38856
rect 67173 38798 70000 38800
rect 67173 38795 67239 38798
rect 69200 38708 70000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 65648 38656 65968 38657
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 38591 65968 38592
rect 0 38028 800 38268
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 50288 38112 50608 38113
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 38047 50608 38048
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 65648 37568 65968 37569
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 37503 65968 37504
rect 66161 37498 66227 37501
rect 69200 37498 70000 37588
rect 66161 37496 70000 37498
rect 66161 37440 66166 37496
rect 66222 37440 70000 37496
rect 66161 37438 70000 37440
rect 66161 37435 66227 37438
rect 69200 37348 70000 37438
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 0 36668 800 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 65648 36480 65968 36481
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 36415 65968 36416
rect 69200 35988 70000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 0 35458 800 35548
rect 4061 35458 4127 35461
rect 0 35456 4127 35458
rect 0 35400 4066 35456
rect 4122 35400 4127 35456
rect 0 35398 4127 35400
rect 0 35308 800 35398
rect 4061 35395 4127 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 65648 35392 65968 35393
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 35327 65968 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 69200 34628 70000 34868
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 65648 34304 65968 34305
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 34239 65968 34240
rect 0 34098 800 34188
rect 3417 34098 3483 34101
rect 0 34096 3483 34098
rect 0 34040 3422 34096
rect 3478 34040 3483 34096
rect 0 34038 3483 34040
rect 0 33948 800 34038
rect 3417 34035 3483 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 66161 33418 66227 33421
rect 69200 33418 70000 33508
rect 66161 33416 70000 33418
rect 66161 33360 66166 33416
rect 66222 33360 70000 33416
rect 66161 33358 70000 33360
rect 66161 33355 66227 33358
rect 69200 33268 70000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 65648 33216 65968 33217
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 33151 65968 33152
rect 0 32588 800 32828
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 65648 32128 65968 32129
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 32063 65968 32064
rect 66069 32058 66135 32061
rect 69200 32058 70000 32148
rect 66069 32056 70000 32058
rect 66069 32000 66074 32056
rect 66130 32000 70000 32056
rect 66069 31998 70000 32000
rect 66069 31995 66135 31998
rect 69200 31908 70000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 0 31378 800 31468
rect 2957 31378 3023 31381
rect 0 31376 3023 31378
rect 0 31320 2962 31376
rect 3018 31320 3023 31376
rect 0 31318 3023 31320
rect 0 31228 800 31318
rect 2957 31315 3023 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 65648 31040 65968 31041
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 30975 65968 30976
rect 66161 30698 66227 30701
rect 69200 30698 70000 30788
rect 66161 30696 70000 30698
rect 66161 30640 66166 30696
rect 66222 30640 70000 30696
rect 66161 30638 70000 30640
rect 66161 30635 66227 30638
rect 69200 30548 70000 30638
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 0 29868 800 30108
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 65648 29952 65968 29953
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 29887 65968 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 69200 29188 70000 29428
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 65648 28864 65968 28865
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 28799 65968 28800
rect 0 28658 800 28748
rect 3417 28658 3483 28661
rect 0 28656 3483 28658
rect 0 28600 3422 28656
rect 3478 28600 3483 28656
rect 0 28598 3483 28600
rect 0 28508 800 28598
rect 3417 28595 3483 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 66161 27978 66227 27981
rect 69200 27978 70000 28068
rect 66161 27976 70000 27978
rect 66161 27920 66166 27976
rect 66222 27920 70000 27976
rect 66161 27918 70000 27920
rect 66161 27915 66227 27918
rect 69200 27828 70000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 65648 27776 65968 27777
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 27711 65968 27712
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 65648 26688 65968 26689
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 26623 65968 26624
rect 66161 26618 66227 26621
rect 69200 26618 70000 26708
rect 66161 26616 70000 26618
rect 66161 26560 66166 26616
rect 66222 26560 70000 26616
rect 66161 26558 70000 26560
rect 66161 26555 66227 26558
rect 69200 26468 70000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 0 25938 800 26028
rect 3141 25938 3207 25941
rect 0 25936 3207 25938
rect 0 25880 3146 25936
rect 3202 25880 3207 25936
rect 0 25878 3207 25880
rect 0 25788 800 25878
rect 3141 25875 3207 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 65648 25600 65968 25601
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 25535 65968 25536
rect 64965 25258 65031 25261
rect 69200 25258 70000 25348
rect 64965 25256 70000 25258
rect 64965 25200 64970 25256
rect 65026 25200 70000 25256
rect 64965 25198 70000 25200
rect 64965 25195 65031 25198
rect 69200 25108 70000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 0 24578 800 24668
rect 3417 24578 3483 24581
rect 0 24576 3483 24578
rect 0 24520 3422 24576
rect 3478 24520 3483 24576
rect 0 24518 3483 24520
rect 0 24428 800 24518
rect 3417 24515 3483 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 65648 24512 65968 24513
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 24447 65968 24448
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 69200 23748 70000 23988
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 65648 23424 65968 23425
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 23359 65968 23360
rect 0 23068 800 23308
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 65648 22336 65968 22337
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 22271 65968 22272
rect 0 21858 800 21948
rect 4061 21858 4127 21861
rect 0 21856 4127 21858
rect 0 21800 4066 21856
rect 4122 21800 4127 21856
rect 0 21798 4127 21800
rect 0 21708 800 21798
rect 4061 21795 4127 21798
rect 66161 21858 66227 21861
rect 69200 21858 70000 21948
rect 66161 21856 70000 21858
rect 66161 21800 66166 21856
rect 66222 21800 70000 21856
rect 66161 21798 70000 21800
rect 66161 21795 66227 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 69200 21708 70000 21798
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 65648 21248 65968 21249
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 21183 65968 21184
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 0 20498 800 20588
rect 4061 20498 4127 20501
rect 0 20496 4127 20498
rect 0 20440 4066 20496
rect 4122 20440 4127 20496
rect 0 20438 4127 20440
rect 0 20348 800 20438
rect 4061 20435 4127 20438
rect 64873 20498 64939 20501
rect 69200 20498 70000 20588
rect 64873 20496 70000 20498
rect 64873 20440 64878 20496
rect 64934 20440 70000 20496
rect 64873 20438 70000 20440
rect 64873 20435 64939 20438
rect 69200 20348 70000 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 65648 20160 65968 20161
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 20095 65968 20096
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 0 18988 800 19228
rect 66161 19138 66227 19141
rect 69200 19138 70000 19228
rect 66161 19136 70000 19138
rect 66161 19080 66166 19136
rect 66222 19080 70000 19136
rect 66161 19078 70000 19080
rect 66161 19075 66227 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 65648 19072 65968 19073
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 19007 65968 19008
rect 69200 18988 70000 19078
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 65648 17984 65968 17985
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 17919 65968 17920
rect 0 17628 800 17868
rect 66161 17778 66227 17781
rect 69200 17778 70000 17868
rect 66161 17776 70000 17778
rect 66161 17720 66166 17776
rect 66222 17720 70000 17776
rect 66161 17718 70000 17720
rect 66161 17715 66227 17718
rect 69200 17628 70000 17718
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 65648 16896 65968 16897
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 16831 65968 16832
rect 0 16418 800 16508
rect 4061 16418 4127 16421
rect 0 16416 4127 16418
rect 0 16360 4066 16416
rect 4122 16360 4127 16416
rect 0 16358 4127 16360
rect 0 16268 800 16358
rect 4061 16355 4127 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 16287 50608 16288
rect 69200 16268 70000 16508
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 65648 15808 65968 15809
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 15743 65968 15744
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 0 15058 800 15148
rect 3969 15058 4035 15061
rect 0 15056 4035 15058
rect 0 15000 3974 15056
rect 4030 15000 4035 15056
rect 0 14998 4035 15000
rect 0 14908 800 14998
rect 3969 14995 4035 14998
rect 69200 14908 70000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 65648 14720 65968 14721
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 14655 65968 14656
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 0 13698 800 13788
rect 4061 13698 4127 13701
rect 0 13696 4127 13698
rect 0 13640 4066 13696
rect 4122 13640 4127 13696
rect 0 13638 4127 13640
rect 0 13548 800 13638
rect 4061 13635 4127 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 65648 13632 65968 13633
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 13567 65968 13568
rect 69200 13548 70000 13788
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 65648 12544 65968 12545
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 12479 65968 12480
rect 0 12188 800 12428
rect 69200 12188 70000 12428
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 65648 11456 65968 11457
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 11391 65968 11392
rect 0 10978 800 11068
rect 3417 10978 3483 10981
rect 0 10976 3483 10978
rect 0 10920 3422 10976
rect 3478 10920 3483 10976
rect 0 10918 3483 10920
rect 0 10828 800 10918
rect 3417 10915 3483 10918
rect 66161 10978 66227 10981
rect 69200 10978 70000 11068
rect 66161 10976 70000 10978
rect 66161 10920 66166 10976
rect 66222 10920 70000 10976
rect 66161 10918 70000 10920
rect 66161 10915 66227 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 69200 10828 70000 10918
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 65648 10368 65968 10369
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 10303 65968 10304
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 0 9618 800 9708
rect 3417 9618 3483 9621
rect 0 9616 3483 9618
rect 0 9560 3422 9616
rect 3478 9560 3483 9616
rect 0 9558 3483 9560
rect 0 9468 800 9558
rect 3417 9555 3483 9558
rect 69200 9468 70000 9708
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 65648 9280 65968 9281
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 9215 65968 9216
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 0 8258 800 8348
rect 3417 8258 3483 8261
rect 0 8256 3483 8258
rect 0 8200 3422 8256
rect 3478 8200 3483 8256
rect 0 8198 3483 8200
rect 0 8108 800 8198
rect 3417 8195 3483 8198
rect 66161 8258 66227 8261
rect 69200 8258 70000 8348
rect 66161 8256 70000 8258
rect 66161 8200 66166 8256
rect 66222 8200 70000 8256
rect 66161 8198 70000 8200
rect 66161 8195 66227 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 65648 8192 65968 8193
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 8127 65968 8128
rect 69200 8108 70000 8198
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 65648 7104 65968 7105
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 7039 65968 7040
rect 0 6898 800 6988
rect 3417 6898 3483 6901
rect 0 6896 3483 6898
rect 0 6840 3422 6896
rect 3478 6840 3483 6896
rect 0 6838 3483 6840
rect 0 6748 800 6838
rect 3417 6835 3483 6838
rect 69200 6748 70000 6988
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 65648 6016 65968 6017
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5951 65968 5952
rect 0 5538 800 5628
rect 3417 5538 3483 5541
rect 0 5536 3483 5538
rect 0 5480 3422 5536
rect 3478 5480 3483 5536
rect 0 5478 3483 5480
rect 0 5388 800 5478
rect 3417 5475 3483 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 69200 5388 70000 5628
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 65648 4928 65968 4929
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 4863 65968 4864
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 0 4178 800 4268
rect 3141 4178 3207 4181
rect 0 4176 3207 4178
rect 0 4120 3146 4176
rect 3202 4120 3207 4176
rect 0 4118 3207 4120
rect 0 4028 800 4118
rect 3141 4115 3207 4118
rect 64781 4178 64847 4181
rect 69200 4178 70000 4268
rect 64781 4176 70000 4178
rect 64781 4120 64786 4176
rect 64842 4120 70000 4176
rect 64781 4118 70000 4120
rect 64781 4115 64847 4118
rect 69200 4028 70000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 65648 3840 65968 3841
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 3775 65968 3776
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 0 2818 800 2908
rect 3509 2818 3575 2821
rect 0 2816 3575 2818
rect 0 2760 3514 2816
rect 3570 2760 3575 2816
rect 0 2758 3575 2760
rect 0 2668 800 2758
rect 3509 2755 3575 2758
rect 66161 2818 66227 2821
rect 69200 2818 70000 2908
rect 66161 2816 70000 2818
rect 66161 2760 66166 2816
rect 66222 2760 70000 2816
rect 66161 2758 70000 2760
rect 66161 2755 66227 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 65648 2752 65968 2753
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2687 65968 2688
rect 69200 2668 70000 2758
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
rect 0 1308 800 1548
rect 65517 1458 65583 1461
rect 69200 1458 70000 1548
rect 65517 1456 70000 1458
rect 65517 1400 65522 1456
rect 65578 1400 70000 1456
rect 65517 1398 70000 1400
rect 65517 1395 65583 1398
rect 69200 1308 70000 1398
rect 69200 -52 70000 188
<< via3 >>
rect 19576 69660 19640 69664
rect 19576 69604 19580 69660
rect 19580 69604 19636 69660
rect 19636 69604 19640 69660
rect 19576 69600 19640 69604
rect 19656 69660 19720 69664
rect 19656 69604 19660 69660
rect 19660 69604 19716 69660
rect 19716 69604 19720 69660
rect 19656 69600 19720 69604
rect 19736 69660 19800 69664
rect 19736 69604 19740 69660
rect 19740 69604 19796 69660
rect 19796 69604 19800 69660
rect 19736 69600 19800 69604
rect 19816 69660 19880 69664
rect 19816 69604 19820 69660
rect 19820 69604 19876 69660
rect 19876 69604 19880 69660
rect 19816 69600 19880 69604
rect 50296 69660 50360 69664
rect 50296 69604 50300 69660
rect 50300 69604 50356 69660
rect 50356 69604 50360 69660
rect 50296 69600 50360 69604
rect 50376 69660 50440 69664
rect 50376 69604 50380 69660
rect 50380 69604 50436 69660
rect 50436 69604 50440 69660
rect 50376 69600 50440 69604
rect 50456 69660 50520 69664
rect 50456 69604 50460 69660
rect 50460 69604 50516 69660
rect 50516 69604 50520 69660
rect 50456 69600 50520 69604
rect 50536 69660 50600 69664
rect 50536 69604 50540 69660
rect 50540 69604 50596 69660
rect 50596 69604 50600 69660
rect 50536 69600 50600 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 34936 69116 35000 69120
rect 34936 69060 34940 69116
rect 34940 69060 34996 69116
rect 34996 69060 35000 69116
rect 34936 69056 35000 69060
rect 35016 69116 35080 69120
rect 35016 69060 35020 69116
rect 35020 69060 35076 69116
rect 35076 69060 35080 69116
rect 35016 69056 35080 69060
rect 35096 69116 35160 69120
rect 35096 69060 35100 69116
rect 35100 69060 35156 69116
rect 35156 69060 35160 69116
rect 35096 69056 35160 69060
rect 35176 69116 35240 69120
rect 35176 69060 35180 69116
rect 35180 69060 35236 69116
rect 35236 69060 35240 69116
rect 35176 69056 35240 69060
rect 65656 69116 65720 69120
rect 65656 69060 65660 69116
rect 65660 69060 65716 69116
rect 65716 69060 65720 69116
rect 65656 69056 65720 69060
rect 65736 69116 65800 69120
rect 65736 69060 65740 69116
rect 65740 69060 65796 69116
rect 65796 69060 65800 69116
rect 65736 69056 65800 69060
rect 65816 69116 65880 69120
rect 65816 69060 65820 69116
rect 65820 69060 65876 69116
rect 65876 69060 65880 69116
rect 65816 69056 65880 69060
rect 65896 69116 65960 69120
rect 65896 69060 65900 69116
rect 65900 69060 65956 69116
rect 65956 69060 65960 69116
rect 65896 69056 65960 69060
rect 19576 68572 19640 68576
rect 19576 68516 19580 68572
rect 19580 68516 19636 68572
rect 19636 68516 19640 68572
rect 19576 68512 19640 68516
rect 19656 68572 19720 68576
rect 19656 68516 19660 68572
rect 19660 68516 19716 68572
rect 19716 68516 19720 68572
rect 19656 68512 19720 68516
rect 19736 68572 19800 68576
rect 19736 68516 19740 68572
rect 19740 68516 19796 68572
rect 19796 68516 19800 68572
rect 19736 68512 19800 68516
rect 19816 68572 19880 68576
rect 19816 68516 19820 68572
rect 19820 68516 19876 68572
rect 19876 68516 19880 68572
rect 19816 68512 19880 68516
rect 50296 68572 50360 68576
rect 50296 68516 50300 68572
rect 50300 68516 50356 68572
rect 50356 68516 50360 68572
rect 50296 68512 50360 68516
rect 50376 68572 50440 68576
rect 50376 68516 50380 68572
rect 50380 68516 50436 68572
rect 50436 68516 50440 68572
rect 50376 68512 50440 68516
rect 50456 68572 50520 68576
rect 50456 68516 50460 68572
rect 50460 68516 50516 68572
rect 50516 68516 50520 68572
rect 50456 68512 50520 68516
rect 50536 68572 50600 68576
rect 50536 68516 50540 68572
rect 50540 68516 50596 68572
rect 50596 68516 50600 68572
rect 50536 68512 50600 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 34936 68028 35000 68032
rect 34936 67972 34940 68028
rect 34940 67972 34996 68028
rect 34996 67972 35000 68028
rect 34936 67968 35000 67972
rect 35016 68028 35080 68032
rect 35016 67972 35020 68028
rect 35020 67972 35076 68028
rect 35076 67972 35080 68028
rect 35016 67968 35080 67972
rect 35096 68028 35160 68032
rect 35096 67972 35100 68028
rect 35100 67972 35156 68028
rect 35156 67972 35160 68028
rect 35096 67968 35160 67972
rect 35176 68028 35240 68032
rect 35176 67972 35180 68028
rect 35180 67972 35236 68028
rect 35236 67972 35240 68028
rect 35176 67968 35240 67972
rect 65656 68028 65720 68032
rect 65656 67972 65660 68028
rect 65660 67972 65716 68028
rect 65716 67972 65720 68028
rect 65656 67968 65720 67972
rect 65736 68028 65800 68032
rect 65736 67972 65740 68028
rect 65740 67972 65796 68028
rect 65796 67972 65800 68028
rect 65736 67968 65800 67972
rect 65816 68028 65880 68032
rect 65816 67972 65820 68028
rect 65820 67972 65876 68028
rect 65876 67972 65880 68028
rect 65816 67968 65880 67972
rect 65896 68028 65960 68032
rect 65896 67972 65900 68028
rect 65900 67972 65956 68028
rect 65956 67972 65960 68028
rect 65896 67968 65960 67972
rect 19576 67484 19640 67488
rect 19576 67428 19580 67484
rect 19580 67428 19636 67484
rect 19636 67428 19640 67484
rect 19576 67424 19640 67428
rect 19656 67484 19720 67488
rect 19656 67428 19660 67484
rect 19660 67428 19716 67484
rect 19716 67428 19720 67484
rect 19656 67424 19720 67428
rect 19736 67484 19800 67488
rect 19736 67428 19740 67484
rect 19740 67428 19796 67484
rect 19796 67428 19800 67484
rect 19736 67424 19800 67428
rect 19816 67484 19880 67488
rect 19816 67428 19820 67484
rect 19820 67428 19876 67484
rect 19876 67428 19880 67484
rect 19816 67424 19880 67428
rect 50296 67484 50360 67488
rect 50296 67428 50300 67484
rect 50300 67428 50356 67484
rect 50356 67428 50360 67484
rect 50296 67424 50360 67428
rect 50376 67484 50440 67488
rect 50376 67428 50380 67484
rect 50380 67428 50436 67484
rect 50436 67428 50440 67484
rect 50376 67424 50440 67428
rect 50456 67484 50520 67488
rect 50456 67428 50460 67484
rect 50460 67428 50516 67484
rect 50516 67428 50520 67484
rect 50456 67424 50520 67428
rect 50536 67484 50600 67488
rect 50536 67428 50540 67484
rect 50540 67428 50596 67484
rect 50596 67428 50600 67484
rect 50536 67424 50600 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 19576 66396 19640 66400
rect 19576 66340 19580 66396
rect 19580 66340 19636 66396
rect 19636 66340 19640 66396
rect 19576 66336 19640 66340
rect 19656 66396 19720 66400
rect 19656 66340 19660 66396
rect 19660 66340 19716 66396
rect 19716 66340 19720 66396
rect 19656 66336 19720 66340
rect 19736 66396 19800 66400
rect 19736 66340 19740 66396
rect 19740 66340 19796 66396
rect 19796 66340 19800 66396
rect 19736 66336 19800 66340
rect 19816 66396 19880 66400
rect 19816 66340 19820 66396
rect 19820 66340 19876 66396
rect 19876 66340 19880 66396
rect 19816 66336 19880 66340
rect 50296 66396 50360 66400
rect 50296 66340 50300 66396
rect 50300 66340 50356 66396
rect 50356 66340 50360 66396
rect 50296 66336 50360 66340
rect 50376 66396 50440 66400
rect 50376 66340 50380 66396
rect 50380 66340 50436 66396
rect 50436 66340 50440 66396
rect 50376 66336 50440 66340
rect 50456 66396 50520 66400
rect 50456 66340 50460 66396
rect 50460 66340 50516 66396
rect 50516 66340 50520 66396
rect 50456 66336 50520 66340
rect 50536 66396 50600 66400
rect 50536 66340 50540 66396
rect 50540 66340 50596 66396
rect 50596 66340 50600 66396
rect 50536 66336 50600 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 19576 65308 19640 65312
rect 19576 65252 19580 65308
rect 19580 65252 19636 65308
rect 19636 65252 19640 65308
rect 19576 65248 19640 65252
rect 19656 65308 19720 65312
rect 19656 65252 19660 65308
rect 19660 65252 19716 65308
rect 19716 65252 19720 65308
rect 19656 65248 19720 65252
rect 19736 65308 19800 65312
rect 19736 65252 19740 65308
rect 19740 65252 19796 65308
rect 19796 65252 19800 65308
rect 19736 65248 19800 65252
rect 19816 65308 19880 65312
rect 19816 65252 19820 65308
rect 19820 65252 19876 65308
rect 19876 65252 19880 65308
rect 19816 65248 19880 65252
rect 50296 65308 50360 65312
rect 50296 65252 50300 65308
rect 50300 65252 50356 65308
rect 50356 65252 50360 65308
rect 50296 65248 50360 65252
rect 50376 65308 50440 65312
rect 50376 65252 50380 65308
rect 50380 65252 50436 65308
rect 50436 65252 50440 65308
rect 50376 65248 50440 65252
rect 50456 65308 50520 65312
rect 50456 65252 50460 65308
rect 50460 65252 50516 65308
rect 50516 65252 50520 65308
rect 50456 65248 50520 65252
rect 50536 65308 50600 65312
rect 50536 65252 50540 65308
rect 50540 65252 50596 65308
rect 50596 65252 50600 65308
rect 50536 65248 50600 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 34936 64764 35000 64768
rect 34936 64708 34940 64764
rect 34940 64708 34996 64764
rect 34996 64708 35000 64764
rect 34936 64704 35000 64708
rect 35016 64764 35080 64768
rect 35016 64708 35020 64764
rect 35020 64708 35076 64764
rect 35076 64708 35080 64764
rect 35016 64704 35080 64708
rect 35096 64764 35160 64768
rect 35096 64708 35100 64764
rect 35100 64708 35156 64764
rect 35156 64708 35160 64764
rect 35096 64704 35160 64708
rect 35176 64764 35240 64768
rect 35176 64708 35180 64764
rect 35180 64708 35236 64764
rect 35236 64708 35240 64764
rect 35176 64704 35240 64708
rect 65656 64764 65720 64768
rect 65656 64708 65660 64764
rect 65660 64708 65716 64764
rect 65716 64708 65720 64764
rect 65656 64704 65720 64708
rect 65736 64764 65800 64768
rect 65736 64708 65740 64764
rect 65740 64708 65796 64764
rect 65796 64708 65800 64764
rect 65736 64704 65800 64708
rect 65816 64764 65880 64768
rect 65816 64708 65820 64764
rect 65820 64708 65876 64764
rect 65876 64708 65880 64764
rect 65816 64704 65880 64708
rect 65896 64764 65960 64768
rect 65896 64708 65900 64764
rect 65900 64708 65956 64764
rect 65956 64708 65960 64764
rect 65896 64704 65960 64708
rect 19576 64220 19640 64224
rect 19576 64164 19580 64220
rect 19580 64164 19636 64220
rect 19636 64164 19640 64220
rect 19576 64160 19640 64164
rect 19656 64220 19720 64224
rect 19656 64164 19660 64220
rect 19660 64164 19716 64220
rect 19716 64164 19720 64220
rect 19656 64160 19720 64164
rect 19736 64220 19800 64224
rect 19736 64164 19740 64220
rect 19740 64164 19796 64220
rect 19796 64164 19800 64220
rect 19736 64160 19800 64164
rect 19816 64220 19880 64224
rect 19816 64164 19820 64220
rect 19820 64164 19876 64220
rect 19876 64164 19880 64220
rect 19816 64160 19880 64164
rect 50296 64220 50360 64224
rect 50296 64164 50300 64220
rect 50300 64164 50356 64220
rect 50356 64164 50360 64220
rect 50296 64160 50360 64164
rect 50376 64220 50440 64224
rect 50376 64164 50380 64220
rect 50380 64164 50436 64220
rect 50436 64164 50440 64220
rect 50376 64160 50440 64164
rect 50456 64220 50520 64224
rect 50456 64164 50460 64220
rect 50460 64164 50516 64220
rect 50516 64164 50520 64220
rect 50456 64160 50520 64164
rect 50536 64220 50600 64224
rect 50536 64164 50540 64220
rect 50540 64164 50596 64220
rect 50596 64164 50600 64220
rect 50536 64160 50600 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 34936 63676 35000 63680
rect 34936 63620 34940 63676
rect 34940 63620 34996 63676
rect 34996 63620 35000 63676
rect 34936 63616 35000 63620
rect 35016 63676 35080 63680
rect 35016 63620 35020 63676
rect 35020 63620 35076 63676
rect 35076 63620 35080 63676
rect 35016 63616 35080 63620
rect 35096 63676 35160 63680
rect 35096 63620 35100 63676
rect 35100 63620 35156 63676
rect 35156 63620 35160 63676
rect 35096 63616 35160 63620
rect 35176 63676 35240 63680
rect 35176 63620 35180 63676
rect 35180 63620 35236 63676
rect 35236 63620 35240 63676
rect 35176 63616 35240 63620
rect 65656 63676 65720 63680
rect 65656 63620 65660 63676
rect 65660 63620 65716 63676
rect 65716 63620 65720 63676
rect 65656 63616 65720 63620
rect 65736 63676 65800 63680
rect 65736 63620 65740 63676
rect 65740 63620 65796 63676
rect 65796 63620 65800 63676
rect 65736 63616 65800 63620
rect 65816 63676 65880 63680
rect 65816 63620 65820 63676
rect 65820 63620 65876 63676
rect 65876 63620 65880 63676
rect 65816 63616 65880 63620
rect 65896 63676 65960 63680
rect 65896 63620 65900 63676
rect 65900 63620 65956 63676
rect 65956 63620 65960 63676
rect 65896 63616 65960 63620
rect 19576 63132 19640 63136
rect 19576 63076 19580 63132
rect 19580 63076 19636 63132
rect 19636 63076 19640 63132
rect 19576 63072 19640 63076
rect 19656 63132 19720 63136
rect 19656 63076 19660 63132
rect 19660 63076 19716 63132
rect 19716 63076 19720 63132
rect 19656 63072 19720 63076
rect 19736 63132 19800 63136
rect 19736 63076 19740 63132
rect 19740 63076 19796 63132
rect 19796 63076 19800 63132
rect 19736 63072 19800 63076
rect 19816 63132 19880 63136
rect 19816 63076 19820 63132
rect 19820 63076 19876 63132
rect 19876 63076 19880 63132
rect 19816 63072 19880 63076
rect 50296 63132 50360 63136
rect 50296 63076 50300 63132
rect 50300 63076 50356 63132
rect 50356 63076 50360 63132
rect 50296 63072 50360 63076
rect 50376 63132 50440 63136
rect 50376 63076 50380 63132
rect 50380 63076 50436 63132
rect 50436 63076 50440 63132
rect 50376 63072 50440 63076
rect 50456 63132 50520 63136
rect 50456 63076 50460 63132
rect 50460 63076 50516 63132
rect 50516 63076 50520 63132
rect 50456 63072 50520 63076
rect 50536 63132 50600 63136
rect 50536 63076 50540 63132
rect 50540 63076 50596 63132
rect 50596 63076 50600 63132
rect 50536 63072 50600 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 34936 62588 35000 62592
rect 34936 62532 34940 62588
rect 34940 62532 34996 62588
rect 34996 62532 35000 62588
rect 34936 62528 35000 62532
rect 35016 62588 35080 62592
rect 35016 62532 35020 62588
rect 35020 62532 35076 62588
rect 35076 62532 35080 62588
rect 35016 62528 35080 62532
rect 35096 62588 35160 62592
rect 35096 62532 35100 62588
rect 35100 62532 35156 62588
rect 35156 62532 35160 62588
rect 35096 62528 35160 62532
rect 35176 62588 35240 62592
rect 35176 62532 35180 62588
rect 35180 62532 35236 62588
rect 35236 62532 35240 62588
rect 35176 62528 35240 62532
rect 65656 62588 65720 62592
rect 65656 62532 65660 62588
rect 65660 62532 65716 62588
rect 65716 62532 65720 62588
rect 65656 62528 65720 62532
rect 65736 62588 65800 62592
rect 65736 62532 65740 62588
rect 65740 62532 65796 62588
rect 65796 62532 65800 62588
rect 65736 62528 65800 62532
rect 65816 62588 65880 62592
rect 65816 62532 65820 62588
rect 65820 62532 65876 62588
rect 65876 62532 65880 62588
rect 65816 62528 65880 62532
rect 65896 62588 65960 62592
rect 65896 62532 65900 62588
rect 65900 62532 65956 62588
rect 65956 62532 65960 62588
rect 65896 62528 65960 62532
rect 19576 62044 19640 62048
rect 19576 61988 19580 62044
rect 19580 61988 19636 62044
rect 19636 61988 19640 62044
rect 19576 61984 19640 61988
rect 19656 62044 19720 62048
rect 19656 61988 19660 62044
rect 19660 61988 19716 62044
rect 19716 61988 19720 62044
rect 19656 61984 19720 61988
rect 19736 62044 19800 62048
rect 19736 61988 19740 62044
rect 19740 61988 19796 62044
rect 19796 61988 19800 62044
rect 19736 61984 19800 61988
rect 19816 62044 19880 62048
rect 19816 61988 19820 62044
rect 19820 61988 19876 62044
rect 19876 61988 19880 62044
rect 19816 61984 19880 61988
rect 50296 62044 50360 62048
rect 50296 61988 50300 62044
rect 50300 61988 50356 62044
rect 50356 61988 50360 62044
rect 50296 61984 50360 61988
rect 50376 62044 50440 62048
rect 50376 61988 50380 62044
rect 50380 61988 50436 62044
rect 50436 61988 50440 62044
rect 50376 61984 50440 61988
rect 50456 62044 50520 62048
rect 50456 61988 50460 62044
rect 50460 61988 50516 62044
rect 50516 61988 50520 62044
rect 50456 61984 50520 61988
rect 50536 62044 50600 62048
rect 50536 61988 50540 62044
rect 50540 61988 50596 62044
rect 50596 61988 50600 62044
rect 50536 61984 50600 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 65656 61500 65720 61504
rect 65656 61444 65660 61500
rect 65660 61444 65716 61500
rect 65716 61444 65720 61500
rect 65656 61440 65720 61444
rect 65736 61500 65800 61504
rect 65736 61444 65740 61500
rect 65740 61444 65796 61500
rect 65796 61444 65800 61500
rect 65736 61440 65800 61444
rect 65816 61500 65880 61504
rect 65816 61444 65820 61500
rect 65820 61444 65876 61500
rect 65876 61444 65880 61500
rect 65816 61440 65880 61444
rect 65896 61500 65960 61504
rect 65896 61444 65900 61500
rect 65900 61444 65956 61500
rect 65956 61444 65960 61500
rect 65896 61440 65960 61444
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 65656 60412 65720 60416
rect 65656 60356 65660 60412
rect 65660 60356 65716 60412
rect 65716 60356 65720 60412
rect 65656 60352 65720 60356
rect 65736 60412 65800 60416
rect 65736 60356 65740 60412
rect 65740 60356 65796 60412
rect 65796 60356 65800 60412
rect 65736 60352 65800 60356
rect 65816 60412 65880 60416
rect 65816 60356 65820 60412
rect 65820 60356 65876 60412
rect 65876 60356 65880 60412
rect 65816 60352 65880 60356
rect 65896 60412 65960 60416
rect 65896 60356 65900 60412
rect 65900 60356 65956 60412
rect 65956 60356 65960 60412
rect 65896 60352 65960 60356
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 65656 59324 65720 59328
rect 65656 59268 65660 59324
rect 65660 59268 65716 59324
rect 65716 59268 65720 59324
rect 65656 59264 65720 59268
rect 65736 59324 65800 59328
rect 65736 59268 65740 59324
rect 65740 59268 65796 59324
rect 65796 59268 65800 59324
rect 65736 59264 65800 59268
rect 65816 59324 65880 59328
rect 65816 59268 65820 59324
rect 65820 59268 65876 59324
rect 65876 59268 65880 59324
rect 65816 59264 65880 59268
rect 65896 59324 65960 59328
rect 65896 59268 65900 59324
rect 65900 59268 65956 59324
rect 65956 59268 65960 59324
rect 65896 59264 65960 59268
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 65656 58236 65720 58240
rect 65656 58180 65660 58236
rect 65660 58180 65716 58236
rect 65716 58180 65720 58236
rect 65656 58176 65720 58180
rect 65736 58236 65800 58240
rect 65736 58180 65740 58236
rect 65740 58180 65796 58236
rect 65796 58180 65800 58236
rect 65736 58176 65800 58180
rect 65816 58236 65880 58240
rect 65816 58180 65820 58236
rect 65820 58180 65876 58236
rect 65876 58180 65880 58236
rect 65816 58176 65880 58180
rect 65896 58236 65960 58240
rect 65896 58180 65900 58236
rect 65900 58180 65956 58236
rect 65956 58180 65960 58236
rect 65896 58176 65960 58180
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 69120 4528 69680
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 65856 4528 66880
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 69664 19888 69680
rect 19568 69600 19576 69664
rect 19640 69600 19656 69664
rect 19720 69600 19736 69664
rect 19800 69600 19816 69664
rect 19880 69600 19888 69664
rect 19568 68576 19888 69600
rect 19568 68512 19576 68576
rect 19640 68512 19656 68576
rect 19720 68512 19736 68576
rect 19800 68512 19816 68576
rect 19880 68512 19888 68576
rect 19568 67488 19888 68512
rect 19568 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19888 67488
rect 19568 66400 19888 67424
rect 19568 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19888 66400
rect 19568 65312 19888 66336
rect 19568 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19888 65312
rect 19568 64224 19888 65248
rect 19568 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19888 64224
rect 19568 63136 19888 64160
rect 19568 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19888 63136
rect 19568 62048 19888 63072
rect 19568 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19888 62048
rect 19568 60960 19888 61984
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 59872 19888 60896
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 69120 35248 69680
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 68032 35248 69056
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 66944 35248 67968
rect 34928 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35248 66944
rect 34928 65856 35248 66880
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 64768 35248 65792
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 63680 35248 64704
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 62592 35248 63616
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 61504 35248 62528
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59328 35248 60352
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 69664 50608 69680
rect 50288 69600 50296 69664
rect 50360 69600 50376 69664
rect 50440 69600 50456 69664
rect 50520 69600 50536 69664
rect 50600 69600 50608 69664
rect 50288 68576 50608 69600
rect 50288 68512 50296 68576
rect 50360 68512 50376 68576
rect 50440 68512 50456 68576
rect 50520 68512 50536 68576
rect 50600 68512 50608 68576
rect 50288 67488 50608 68512
rect 50288 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50608 67488
rect 50288 66400 50608 67424
rect 50288 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50608 66400
rect 50288 65312 50608 66336
rect 50288 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50608 65312
rect 50288 64224 50608 65248
rect 50288 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50608 64224
rect 50288 63136 50608 64160
rect 50288 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50608 63136
rect 50288 62048 50608 63072
rect 50288 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50608 62048
rect 50288 60960 50608 61984
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 69120 65968 69680
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 68032 65968 69056
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 66944 65968 67968
rect 65648 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65968 66944
rect 65648 65856 65968 66880
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 64768 65968 65792
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 63680 65968 64704
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 62592 65968 63616
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 61504 65968 62528
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 60416 65968 61440
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 59328 65968 60352
rect 65648 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65968 59328
rect 65648 58240 65968 59264
rect 65648 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65968 58240
rect 65648 57152 65968 58176
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
use sky130_fd_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1644511149
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1644511149
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_405
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1644511149
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1644511149
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_489
timestamp 1644511149
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1644511149
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_517
timestamp 1644511149
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1644511149
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_545
timestamp 1644511149
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1644511149
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_561
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1644511149
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_589
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_601
timestamp 1644511149
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1644511149
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_617
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_629
timestamp 1644511149
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1644511149
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_645
timestamp 1644511149
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_657
timestamp 1644511149
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1644511149
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_673
timestamp 1644511149
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_685
timestamp 1644511149
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1644511149
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_701
timestamp 1644511149
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_713
timestamp 1644511149
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1644511149
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_417
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_429
timestamp 1644511149
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1644511149
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_461
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_473
timestamp 1644511149
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_485
timestamp 1644511149
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1644511149
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1644511149
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_529
timestamp 1644511149
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_541
timestamp 1644511149
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1644511149
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1644511149
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_573
timestamp 1644511149
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_585
timestamp 1644511149
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_597
timestamp 1644511149
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1644511149
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1644511149
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_617
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_629
timestamp 1644511149
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_641
timestamp 1644511149
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_653
timestamp 1644511149
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1644511149
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1644511149
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_673
timestamp 1644511149
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_685
timestamp 1644511149
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_697
timestamp 1644511149
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_709
timestamp 1644511149
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1644511149
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1644511149
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1644511149
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_330
timestamp 1644511149
transform 1 0 31464 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_342
timestamp 1644511149
transform 1 0 32568 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_354 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_489
timestamp 1644511149
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_501
timestamp 1644511149
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_513
timestamp 1644511149
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1644511149
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1644511149
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_613
timestamp 1644511149
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_625
timestamp 1644511149
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1644511149
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1644511149
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_645
timestamp 1644511149
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_657
timestamp 1644511149
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_669
timestamp 1644511149
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_681
timestamp 1644511149
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1644511149
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1644511149
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_701
timestamp 1644511149
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_713
timestamp 1644511149
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_725
timestamp 1644511149
transform 1 0 67804 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_121
timestamp 1644511149
transform 1 0 12236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_126
timestamp 1644511149
transform 1 0 12696 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_138
timestamp 1644511149
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_150
timestamp 1644511149
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1644511149
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_299
timestamp 1644511149
transform 1 0 28612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_324
timestamp 1644511149
transform 1 0 30912 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_629
timestamp 1644511149
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_641
timestamp 1644511149
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_653
timestamp 1644511149
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1644511149
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1644511149
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_673
timestamp 1644511149
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_685
timestamp 1644511149
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_697
timestamp 1644511149
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_709
timestamp 1644511149
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1644511149
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1644511149
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_729
timestamp 1644511149
transform 1 0 68172 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_312
timestamp 1644511149
transform 1 0 29808 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_324
timestamp 1644511149
transform 1 0 30912 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_336
timestamp 1644511149
transform 1 0 32016 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_348
timestamp 1644511149
transform 1 0 33120 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1644511149
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_625
timestamp 1644511149
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1644511149
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1644511149
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_645
timestamp 1644511149
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_657
timestamp 1644511149
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_669
timestamp 1644511149
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_681
timestamp 1644511149
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1644511149
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1644511149
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_701
timestamp 1644511149
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_713
timestamp 1644511149
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_725
timestamp 1644511149
transform 1 0 67804 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_124
timestamp 1644511149
transform 1 0 12512 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_136
timestamp 1644511149
transform 1 0 13616 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_148
timestamp 1644511149
transform 1 0 14720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 1644511149
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_457
timestamp 1644511149
transform 1 0 43148 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_481
timestamp 1644511149
transform 1 0 45356 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_493
timestamp 1644511149
transform 1 0 46460 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_501
timestamp 1644511149
transform 1 0 47196 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_629
timestamp 1644511149
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_641
timestamp 1644511149
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_653
timestamp 1644511149
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1644511149
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1644511149
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_673
timestamp 1644511149
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_685
timestamp 1644511149
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_697
timestamp 1644511149
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_709
timestamp 1644511149
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1644511149
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1644511149
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_729
timestamp 1644511149
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_130
timestamp 1644511149
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1644511149
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_464
timestamp 1644511149
transform 1 0 43792 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_625
timestamp 1644511149
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1644511149
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1644511149
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_645
timestamp 1644511149
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_657
timestamp 1644511149
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_669
timestamp 1644511149
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_681
timestamp 1644511149
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1644511149
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1644511149
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_701
timestamp 1644511149
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_713
timestamp 1644511149
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_725
timestamp 1644511149
transform 1 0 67804 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1644511149
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_134
timestamp 1644511149
transform 1 0 13432 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_146
timestamp 1644511149
transform 1 0 14536 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_158
timestamp 1644511149
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1644511149
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_457
timestamp 1644511149
transform 1 0 43148 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_462
timestamp 1644511149
transform 1 0 43608 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_474
timestamp 1644511149
transform 1 0 44712 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_486
timestamp 1644511149
transform 1 0 45816 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_498
timestamp 1644511149
transform 1 0 46920 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_629
timestamp 1644511149
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_641
timestamp 1644511149
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_653
timestamp 1644511149
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1644511149
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1644511149
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_673
timestamp 1644511149
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_685
timestamp 1644511149
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_697
timestamp 1644511149
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_709
timestamp 1644511149
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1644511149
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1644511149
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_729
timestamp 1644511149
transform 1 0 68172 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_103
timestamp 1644511149
transform 1 0 10580 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_107
timestamp 1644511149
transform 1 0 10948 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_114
timestamp 1644511149
transform 1 0 11592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_625
timestamp 1644511149
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1644511149
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1644511149
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_645
timestamp 1644511149
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_657
timestamp 1644511149
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_669
timestamp 1644511149
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_681
timestamp 1644511149
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1644511149
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1644511149
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_701
timestamp 1644511149
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_713
timestamp 1644511149
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_725
timestamp 1644511149
transform 1 0 67804 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_629
timestamp 1644511149
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_641
timestamp 1644511149
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_653
timestamp 1644511149
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1644511149
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1644511149
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_673
timestamp 1644511149
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_685
timestamp 1644511149
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_697
timestamp 1644511149
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_709
timestamp 1644511149
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1644511149
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1644511149
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_729
timestamp 1644511149
transform 1 0 68172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_497
timestamp 1644511149
transform 1 0 46828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_503
timestamp 1644511149
transform 1 0 47380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_528
timestamp 1644511149
transform 1 0 49680 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_625
timestamp 1644511149
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1644511149
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1644511149
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_645
timestamp 1644511149
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_657
timestamp 1644511149
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_669
timestamp 1644511149
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_681
timestamp 1644511149
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1644511149
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1644511149
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_701
timestamp 1644511149
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_713
timestamp 1644511149
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_725
timestamp 1644511149
transform 1 0 67804 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_511
timestamp 1644511149
transform 1 0 48116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_523
timestamp 1644511149
transform 1 0 49220 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_535
timestamp 1644511149
transform 1 0 50324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_547
timestamp 1644511149
transform 1 0 51428 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_629
timestamp 1644511149
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_641
timestamp 1644511149
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_653
timestamp 1644511149
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1644511149
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1644511149
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_673
timestamp 1644511149
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_685
timestamp 1644511149
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_697
timestamp 1644511149
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_709
timestamp 1644511149
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1644511149
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1644511149
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_729
timestamp 1644511149
transform 1 0 68172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_625
timestamp 1644511149
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1644511149
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1644511149
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_645
timestamp 1644511149
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_657
timestamp 1644511149
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_669
timestamp 1644511149
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_681
timestamp 1644511149
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1644511149
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1644511149
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_701
timestamp 1644511149
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_713
timestamp 1644511149
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_725
timestamp 1644511149
transform 1 0 67804 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_401
timestamp 1644511149
transform 1 0 37996 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_423
timestamp 1644511149
transform 1 0 40020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_435
timestamp 1644511149
transform 1 0 41124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_629
timestamp 1644511149
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_641
timestamp 1644511149
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_653
timestamp 1644511149
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1644511149
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1644511149
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_673
timestamp 1644511149
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_685
timestamp 1644511149
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_697
timestamp 1644511149
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_709
timestamp 1644511149
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1644511149
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1644511149
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_729
timestamp 1644511149
transform 1 0 68172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1644511149
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_115
timestamp 1644511149
transform 1 0 11684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_127
timestamp 1644511149
transform 1 0 12788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_293
timestamp 1644511149
transform 1 0 28060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1644511149
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_498
timestamp 1644511149
transform 1 0 46920 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_510
timestamp 1644511149
transform 1 0 48024 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_522
timestamp 1644511149
transform 1 0 49128 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_530
timestamp 1644511149
transform 1 0 49864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_625
timestamp 1644511149
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1644511149
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1644511149
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_645
timestamp 1644511149
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_657
timestamp 1644511149
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_669
timestamp 1644511149
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_681
timestamp 1644511149
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1644511149
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1644511149
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_701
timestamp 1644511149
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_713
timestamp 1644511149
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_725
timestamp 1644511149
transform 1 0 67804 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_89
timestamp 1644511149
transform 1 0 9292 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_100
timestamp 1644511149
transform 1 0 10304 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_255
timestamp 1644511149
transform 1 0 24564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_259
timestamp 1644511149
transform 1 0 24932 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_271
timestamp 1644511149
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_308
timestamp 1644511149
transform 1 0 29440 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_320
timestamp 1644511149
transform 1 0 30544 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1644511149
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_401
timestamp 1644511149
transform 1 0 37996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_406
timestamp 1644511149
transform 1 0 38456 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_413
timestamp 1644511149
transform 1 0 39100 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_425
timestamp 1644511149
transform 1 0 40204 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_437
timestamp 1644511149
transform 1 0 41308 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_445
timestamp 1644511149
transform 1 0 42044 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_465
timestamp 1644511149
transform 1 0 43884 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_469
timestamp 1644511149
transform 1 0 44252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_476
timestamp 1644511149
transform 1 0 44896 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_488
timestamp 1644511149
transform 1 0 46000 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_629
timestamp 1644511149
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_641
timestamp 1644511149
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_653
timestamp 1644511149
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1644511149
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1644511149
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_673
timestamp 1644511149
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_685
timestamp 1644511149
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_697
timestamp 1644511149
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_709
timestamp 1644511149
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1644511149
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1644511149
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_729
timestamp 1644511149
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_106
timestamp 1644511149
transform 1 0 10856 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_118
timestamp 1644511149
transform 1 0 11960 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 1644511149
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1644511149
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_274
timestamp 1644511149
transform 1 0 26312 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_286
timestamp 1644511149
transform 1 0 27416 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_290
timestamp 1644511149
transform 1 0 27784 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_302
timestamp 1644511149
transform 1 0 28888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_426
timestamp 1644511149
transform 1 0 40296 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_438
timestamp 1644511149
transform 1 0 41400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_462
timestamp 1644511149
transform 1 0 43608 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1644511149
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_625
timestamp 1644511149
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1644511149
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1644511149
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_645
timestamp 1644511149
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_657
timestamp 1644511149
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_669
timestamp 1644511149
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_681
timestamp 1644511149
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1644511149
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1644511149
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_701
timestamp 1644511149
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_713
timestamp 1644511149
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_725
timestamp 1644511149
transform 1 0 67804 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_77
timestamp 1644511149
transform 1 0 8188 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1644511149
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1644511149
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_254
timestamp 1644511149
transform 1 0 24472 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_266
timestamp 1644511149
transform 1 0 25576 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1644511149
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_444
timestamp 1644511149
transform 1 0 41952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_452
timestamp 1644511149
transform 1 0 42688 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_464
timestamp 1644511149
transform 1 0 43792 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_476
timestamp 1644511149
transform 1 0 44896 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_488
timestamp 1644511149
transform 1 0 46000 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_500
timestamp 1644511149
transform 1 0 47104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_629
timestamp 1644511149
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_641
timestamp 1644511149
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_653
timestamp 1644511149
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1644511149
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1644511149
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_673
timestamp 1644511149
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_685
timestamp 1644511149
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_697
timestamp 1644511149
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_709
timestamp 1644511149
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1644511149
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1644511149
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_729
timestamp 1644511149
transform 1 0 68172 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_73
timestamp 1644511149
transform 1 0 7820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1644511149
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_94
timestamp 1644511149
transform 1 0 9752 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_106
timestamp 1644511149
transform 1 0 10856 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_118
timestamp 1644511149
transform 1 0 11960 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_130
timestamp 1644511149
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1644511149
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_428
timestamp 1644511149
transform 1 0 40480 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_436
timestamp 1644511149
transform 1 0 41216 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_442
timestamp 1644511149
transform 1 0 41768 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_454
timestamp 1644511149
transform 1 0 42872 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_466
timestamp 1644511149
transform 1 0 43976 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_474
timestamp 1644511149
transform 1 0 44712 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_625
timestamp 1644511149
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1644511149
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1644511149
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_645
timestamp 1644511149
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_657
timestamp 1644511149
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_669
timestamp 1644511149
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_681
timestamp 1644511149
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1644511149
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1644511149
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_701
timestamp 1644511149
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_713
timestamp 1644511149
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_725
timestamp 1644511149
transform 1 0 67804 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_85
timestamp 1644511149
transform 1 0 8924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_89
timestamp 1644511149
transform 1 0 9292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_101
timestamp 1644511149
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1644511149
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_116
timestamp 1644511149
transform 1 0 11776 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_128
timestamp 1644511149
transform 1 0 12880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_140
timestamp 1644511149
transform 1 0 13984 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_152
timestamp 1644511149
transform 1 0 15088 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_629
timestamp 1644511149
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_641
timestamp 1644511149
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_653
timestamp 1644511149
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1644511149
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1644511149
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_673
timestamp 1644511149
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_685
timestamp 1644511149
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_697
timestamp 1644511149
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_709
timestamp 1644511149
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1644511149
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1644511149
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_729
timestamp 1644511149
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_122
timestamp 1644511149
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1644511149
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_149
timestamp 1644511149
transform 1 0 14812 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_171
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_183
timestamp 1644511149
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_338
timestamp 1644511149
transform 1 0 32200 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_350
timestamp 1644511149
transform 1 0 33304 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1644511149
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_373
timestamp 1644511149
transform 1 0 35420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_396
timestamp 1644511149
transform 1 0 37536 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_408
timestamp 1644511149
transform 1 0 38640 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_625
timestamp 1644511149
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1644511149
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1644511149
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_645
timestamp 1644511149
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_657
timestamp 1644511149
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_669
timestamp 1644511149
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_681
timestamp 1644511149
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1644511149
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1644511149
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_701
timestamp 1644511149
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_713
timestamp 1644511149
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_725
timestamp 1644511149
transform 1 0 67804 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_101
timestamp 1644511149
transform 1 0 10396 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_154
timestamp 1644511149
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1644511149
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_323
timestamp 1644511149
transform 1 0 30820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 1644511149
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_629
timestamp 1644511149
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_641
timestamp 1644511149
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_653
timestamp 1644511149
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1644511149
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1644511149
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_673
timestamp 1644511149
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_685
timestamp 1644511149
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_697
timestamp 1644511149
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_709
timestamp 1644511149
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1644511149
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1644511149
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_729
timestamp 1644511149
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1644511149
transform 1 0 15272 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1644511149
transform 1 0 16376 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1644511149
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_373
timestamp 1644511149
transform 1 0 35420 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_379
timestamp 1644511149
transform 1 0 35972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_386
timestamp 1644511149
transform 1 0 36616 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_398
timestamp 1644511149
transform 1 0 37720 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_410
timestamp 1644511149
transform 1 0 38824 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1644511149
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_625
timestamp 1644511149
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1644511149
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1644511149
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_645
timestamp 1644511149
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_657
timestamp 1644511149
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_669
timestamp 1644511149
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_681
timestamp 1644511149
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1644511149
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1644511149
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_701
timestamp 1644511149
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_713
timestamp 1644511149
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_725
timestamp 1644511149
transform 1 0 67804 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_260
timestamp 1644511149
transform 1 0 25024 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1644511149
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_629
timestamp 1644511149
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_641
timestamp 1644511149
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_653
timestamp 1644511149
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1644511149
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1644511149
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_694
timestamp 1644511149
transform 1 0 64952 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_706
timestamp 1644511149
transform 1 0 66056 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_718
timestamp 1644511149
transform 1 0 67160 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_726
timestamp 1644511149
transform 1 0 67896 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_729
timestamp 1644511149
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_237
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_241
timestamp 1644511149
transform 1 0 23276 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_625
timestamp 1644511149
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1644511149
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1644511149
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_645
timestamp 1644511149
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_657
timestamp 1644511149
transform 1 0 61548 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_661
timestamp 1644511149
transform 1 0 61916 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_665
timestamp 1644511149
transform 1 0 62284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_672
timestamp 1644511149
transform 1 0 62928 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_684
timestamp 1644511149
transform 1 0 64032 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_696
timestamp 1644511149
transform 1 0 65136 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_701
timestamp 1644511149
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_713
timestamp 1644511149
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_725
timestamp 1644511149
transform 1 0 67804 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_629
timestamp 1644511149
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_641
timestamp 1644511149
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_653
timestamp 1644511149
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1644511149
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1644511149
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_673
timestamp 1644511149
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_685
timestamp 1644511149
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_697
timestamp 1644511149
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_709
timestamp 1644511149
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1644511149
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1644511149
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_729
timestamp 1644511149
transform 1 0 68172 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1644511149
transform 1 0 14352 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1644511149
transform 1 0 15456 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1644511149
transform 1 0 16560 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1644511149
transform 1 0 17664 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_625
timestamp 1644511149
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1644511149
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1644511149
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_645
timestamp 1644511149
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_657
timestamp 1644511149
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_669
timestamp 1644511149
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_681
timestamp 1644511149
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1644511149
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1644511149
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_701
timestamp 1644511149
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_713
timestamp 1644511149
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_725
timestamp 1644511149
transform 1 0 67804 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1644511149
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_396
timestamp 1644511149
transform 1 0 37536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_408
timestamp 1644511149
transform 1 0 38640 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_420
timestamp 1644511149
transform 1 0 39744 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_432
timestamp 1644511149
transform 1 0 40848 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_444
timestamp 1644511149
transform 1 0 41952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_629
timestamp 1644511149
transform 1 0 58972 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_652
timestamp 1644511149
transform 1 0 61088 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_664
timestamp 1644511149
transform 1 0 62192 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_673
timestamp 1644511149
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_685
timestamp 1644511149
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_697
timestamp 1644511149
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_709
timestamp 1644511149
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1644511149
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1644511149
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_729
timestamp 1644511149
transform 1 0 68172 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1644511149
transform 1 0 14352 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1644511149
transform 1 0 15456 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1644511149
transform 1 0 16560 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1644511149
transform 1 0 17664 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_384
timestamp 1644511149
transform 1 0 36432 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_409
timestamp 1644511149
transform 1 0 38732 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_417
timestamp 1644511149
transform 1 0 39468 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_625
timestamp 1644511149
transform 1 0 58604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_630
timestamp 1644511149
transform 1 0 59064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1644511149
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1644511149
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_645
timestamp 1644511149
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_657
timestamp 1644511149
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_669
timestamp 1644511149
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_681
timestamp 1644511149
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1644511149
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1644511149
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_701
timestamp 1644511149
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_713
timestamp 1644511149
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_725
timestamp 1644511149
transform 1 0 67804 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_271
timestamp 1644511149
transform 1 0 26036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_629
timestamp 1644511149
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_641
timestamp 1644511149
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_653
timestamp 1644511149
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1644511149
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1644511149
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_673
timestamp 1644511149
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_685
timestamp 1644511149
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_697
timestamp 1644511149
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_709
timestamp 1644511149
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1644511149
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1644511149
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_729
timestamp 1644511149
transform 1 0 68172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_258
timestamp 1644511149
transform 1 0 24840 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_270
timestamp 1644511149
transform 1 0 25944 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_282
timestamp 1644511149
transform 1 0 27048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_373
timestamp 1644511149
transform 1 0 35420 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_395
timestamp 1644511149
transform 1 0 37444 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_407
timestamp 1644511149
transform 1 0 38548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_625
timestamp 1644511149
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1644511149
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1644511149
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_645
timestamp 1644511149
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_657
timestamp 1644511149
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_669
timestamp 1644511149
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_681
timestamp 1644511149
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1644511149
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1644511149
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_701
timestamp 1644511149
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_713
timestamp 1644511149
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_725
timestamp 1644511149
transform 1 0 67804 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_289
timestamp 1644511149
transform 1 0 27692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_294
timestamp 1644511149
transform 1 0 28152 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_301
timestamp 1644511149
transform 1 0 28796 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_313
timestamp 1644511149
transform 1 0 29900 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_325
timestamp 1644511149
transform 1 0 31004 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1644511149
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_369
timestamp 1644511149
transform 1 0 35052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_380
timestamp 1644511149
transform 1 0 36064 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_629
timestamp 1644511149
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_641
timestamp 1644511149
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_653
timestamp 1644511149
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1644511149
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1644511149
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_673
timestamp 1644511149
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_685
timestamp 1644511149
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_697
timestamp 1644511149
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_709
timestamp 1644511149
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1644511149
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1644511149
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_729
timestamp 1644511149
transform 1 0 68172 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_88
timestamp 1644511149
transform 1 0 9200 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_100
timestamp 1644511149
transform 1 0 10304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_112
timestamp 1644511149
transform 1 0 11408 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_124
timestamp 1644511149
transform 1 0 12512 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_625
timestamp 1644511149
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1644511149
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1644511149
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_645
timestamp 1644511149
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_657
timestamp 1644511149
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_669
timestamp 1644511149
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_681
timestamp 1644511149
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1644511149
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1644511149
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_701
timestamp 1644511149
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_713
timestamp 1644511149
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_725
timestamp 1644511149
transform 1 0 67804 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_103
timestamp 1644511149
transform 1 0 10580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_629
timestamp 1644511149
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_641
timestamp 1644511149
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_653
timestamp 1644511149
transform 1 0 61180 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_661
timestamp 1644511149
transform 1 0 61916 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_667
timestamp 1644511149
transform 1 0 62468 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1644511149
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_694
timestamp 1644511149
transform 1 0 64952 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_706
timestamp 1644511149
transform 1 0 66056 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_718
timestamp 1644511149
transform 1 0 67160 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_726
timestamp 1644511149
transform 1 0 67896 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_729
timestamp 1644511149
transform 1 0 68172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_88
timestamp 1644511149
transform 1 0 9200 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_100
timestamp 1644511149
transform 1 0 10304 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_112
timestamp 1644511149
transform 1 0 11408 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_124
timestamp 1644511149
transform 1 0 12512 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_625
timestamp 1644511149
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1644511149
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1644511149
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_645
timestamp 1644511149
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_657
timestamp 1644511149
transform 1 0 61548 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_665
timestamp 1644511149
transform 1 0 62284 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_670
timestamp 1644511149
transform 1 0 62744 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_682
timestamp 1644511149
transform 1 0 63848 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_694
timestamp 1644511149
transform 1 0 64952 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_701
timestamp 1644511149
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_713
timestamp 1644511149
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_725
timestamp 1644511149
transform 1 0 67804 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_60
timestamp 1644511149
transform 1 0 6624 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_72
timestamp 1644511149
transform 1 0 7728 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_84
timestamp 1644511149
transform 1 0 8832 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_95
timestamp 1644511149
transform 1 0 9844 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp 1644511149
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_117
timestamp 1644511149
transform 1 0 11868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_121
timestamp 1644511149
transform 1 0 12236 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_133
timestamp 1644511149
transform 1 0 13340 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_145
timestamp 1644511149
transform 1 0 14444 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_157
timestamp 1644511149
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1644511149
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_602
timestamp 1644511149
transform 1 0 56488 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_614
timestamp 1644511149
transform 1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_629
timestamp 1644511149
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_641
timestamp 1644511149
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_653
timestamp 1644511149
transform 1 0 61180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_657
timestamp 1644511149
transform 1 0 61548 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_661
timestamp 1644511149
transform 1 0 61916 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_669
timestamp 1644511149
transform 1 0 62652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_673
timestamp 1644511149
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_685
timestamp 1644511149
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_697
timestamp 1644511149
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_709
timestamp 1644511149
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1644511149
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1644511149
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_729
timestamp 1644511149
transform 1 0 68172 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_49
timestamp 1644511149
transform 1 0 5612 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_71
timestamp 1644511149
transform 1 0 7636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1644511149
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_114
timestamp 1644511149
transform 1 0 11592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_268
timestamp 1644511149
transform 1 0 25760 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_293
timestamp 1644511149
transform 1 0 28060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1644511149
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_556
timestamp 1644511149
transform 1 0 52256 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_568
timestamp 1644511149
transform 1 0 53360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_580
timestamp 1644511149
transform 1 0 54464 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_597
timestamp 1644511149
transform 1 0 56028 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_621
timestamp 1644511149
transform 1 0 58236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_633
timestamp 1644511149
transform 1 0 59340 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_641
timestamp 1644511149
transform 1 0 60076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_645
timestamp 1644511149
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_657
timestamp 1644511149
transform 1 0 61548 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_680
timestamp 1644511149
transform 1 0 63664 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_692
timestamp 1644511149
transform 1 0 64768 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_701
timestamp 1644511149
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_713
timestamp 1644511149
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_725
timestamp 1644511149
transform 1 0 67804 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_60
timestamp 1644511149
transform 1 0 6624 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_72
timestamp 1644511149
transform 1 0 7728 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_84
timestamp 1644511149
transform 1 0 8832 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_88
timestamp 1644511149
transform 1 0 9200 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_92
timestamp 1644511149
transform 1 0 9568 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_104
timestamp 1644511149
transform 1 0 10672 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_119
timestamp 1644511149
transform 1 0 12052 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_131
timestamp 1644511149
transform 1 0 13156 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_143
timestamp 1644511149
transform 1 0 14260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_155
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_552
timestamp 1644511149
transform 1 0 51888 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_582
timestamp 1644511149
transform 1 0 54648 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_594
timestamp 1644511149
transform 1 0 55752 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_600
timestamp 1644511149
transform 1 0 56304 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_604
timestamp 1644511149
transform 1 0 56672 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_629
timestamp 1644511149
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_641
timestamp 1644511149
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_653
timestamp 1644511149
transform 1 0 61180 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_659
timestamp 1644511149
transform 1 0 61732 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_663
timestamp 1644511149
transform 1 0 62100 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1644511149
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_673
timestamp 1644511149
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_685
timestamp 1644511149
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_697
timestamp 1644511149
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_709
timestamp 1644511149
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1644511149
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1644511149
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_729
timestamp 1644511149
transform 1 0 68172 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_625
timestamp 1644511149
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1644511149
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1644511149
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_645
timestamp 1644511149
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_657
timestamp 1644511149
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_669
timestamp 1644511149
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_681
timestamp 1644511149
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1644511149
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1644511149
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_701
timestamp 1644511149
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_713
timestamp 1644511149
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_725
timestamp 1644511149
transform 1 0 67804 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_259
timestamp 1644511149
transform 1 0 24932 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_271
timestamp 1644511149
transform 1 0 26036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_629
timestamp 1644511149
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_641
timestamp 1644511149
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_653
timestamp 1644511149
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1644511149
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1644511149
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_673
timestamp 1644511149
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_685
timestamp 1644511149
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_697
timestamp 1644511149
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_709
timestamp 1644511149
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1644511149
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1644511149
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_729
timestamp 1644511149
transform 1 0 68172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_127
timestamp 1644511149
transform 1 0 12788 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_131
timestamp 1644511149
transform 1 0 13156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_300
timestamp 1644511149
transform 1 0 28704 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_625
timestamp 1644511149
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1644511149
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1644511149
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_645
timestamp 1644511149
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_657
timestamp 1644511149
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_669
timestamp 1644511149
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_681
timestamp 1644511149
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1644511149
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1644511149
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_701
timestamp 1644511149
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_713
timestamp 1644511149
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_725
timestamp 1644511149
transform 1 0 67804 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_121
timestamp 1644511149
transform 1 0 12236 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_143
timestamp 1644511149
transform 1 0 14260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_155
timestamp 1644511149
transform 1 0 15364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_233
timestamp 1644511149
transform 1 0 22540 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1644511149
transform 1 0 23092 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_246
timestamp 1644511149
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_258
timestamp 1644511149
transform 1 0 24840 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1644511149
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1644511149
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_315
timestamp 1644511149
transform 1 0 30084 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_358
timestamp 1644511149
transform 1 0 34040 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_370
timestamp 1644511149
transform 1 0 35144 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_382
timestamp 1644511149
transform 1 0 36248 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1644511149
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_629
timestamp 1644511149
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_641
timestamp 1644511149
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_653
timestamp 1644511149
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1644511149
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1644511149
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_673
timestamp 1644511149
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_685
timestamp 1644511149
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_697
timestamp 1644511149
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_709
timestamp 1644511149
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1644511149
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1644511149
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_729
timestamp 1644511149
transform 1 0 68172 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1644511149
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_290
timestamp 1644511149
transform 1 0 27784 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_297
timestamp 1644511149
transform 1 0 28428 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1644511149
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_339
timestamp 1644511149
transform 1 0 32292 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_346
timestamp 1644511149
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_358
timestamp 1644511149
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_625
timestamp 1644511149
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1644511149
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1644511149
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_645
timestamp 1644511149
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_657
timestamp 1644511149
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_669
timestamp 1644511149
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_681
timestamp 1644511149
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1644511149
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1644511149
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_701
timestamp 1644511149
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_713
timestamp 1644511149
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_725
timestamp 1644511149
transform 1 0 67804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_284
timestamp 1644511149
transform 1 0 27232 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_296
timestamp 1644511149
transform 1 0 28336 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_308
timestamp 1644511149
transform 1 0 29440 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_320
timestamp 1644511149
transform 1 0 30544 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_603
timestamp 1644511149
transform 1 0 56580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_623
timestamp 1644511149
transform 1 0 58420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_635
timestamp 1644511149
transform 1 0 59524 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_647
timestamp 1644511149
transform 1 0 60628 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_659
timestamp 1644511149
transform 1 0 61732 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1644511149
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_673
timestamp 1644511149
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_685
timestamp 1644511149
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_697
timestamp 1644511149
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_709
timestamp 1644511149
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1644511149
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1644511149
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_729
timestamp 1644511149
transform 1 0 68172 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_269
timestamp 1644511149
transform 1 0 25852 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_273
timestamp 1644511149
transform 1 0 26220 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_285
timestamp 1644511149
transform 1 0 27324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_297
timestamp 1644511149
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1644511149
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_353
timestamp 1644511149
transform 1 0 33580 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_358
timestamp 1644511149
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_368
timestamp 1644511149
transform 1 0 34960 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_380
timestamp 1644511149
transform 1 0 36064 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_392
timestamp 1644511149
transform 1 0 37168 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_404
timestamp 1644511149
transform 1 0 38272 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1644511149
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_593
timestamp 1644511149
transform 1 0 55660 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_615
timestamp 1644511149
transform 1 0 57684 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_640
timestamp 1644511149
transform 1 0 59984 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_645
timestamp 1644511149
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_657
timestamp 1644511149
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_669
timestamp 1644511149
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_681
timestamp 1644511149
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1644511149
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1644511149
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_701
timestamp 1644511149
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_713
timestamp 1644511149
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_725
timestamp 1644511149
transform 1 0 67804 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_376
timestamp 1644511149
transform 1 0 35696 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1644511149
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_604
timestamp 1644511149
transform 1 0 56672 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_624
timestamp 1644511149
transform 1 0 58512 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_636
timestamp 1644511149
transform 1 0 59616 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_648
timestamp 1644511149
transform 1 0 60720 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_660
timestamp 1644511149
transform 1 0 61824 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_673
timestamp 1644511149
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_685
timestamp 1644511149
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_697
timestamp 1644511149
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_709
timestamp 1644511149
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1644511149
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1644511149
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_729
timestamp 1644511149
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_539
timestamp 1644511149
transform 1 0 50692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_551
timestamp 1644511149
transform 1 0 51796 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_563
timestamp 1644511149
transform 1 0 52900 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_575
timestamp 1644511149
transform 1 0 54004 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1644511149
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_613
timestamp 1644511149
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_625
timestamp 1644511149
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1644511149
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1644511149
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_645
timestamp 1644511149
transform 1 0 60444 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_651
timestamp 1644511149
transform 1 0 60996 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_655
timestamp 1644511149
transform 1 0 61364 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_667
timestamp 1644511149
transform 1 0 62468 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_679
timestamp 1644511149
transform 1 0 63572 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_691
timestamp 1644511149
transform 1 0 64676 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1644511149
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_701
timestamp 1644511149
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_713
timestamp 1644511149
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_725
timestamp 1644511149
transform 1 0 67804 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_525
timestamp 1644511149
transform 1 0 49404 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_531
timestamp 1644511149
transform 1 0 49956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_556
timestamp 1644511149
transform 1 0 52256 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1644511149
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_629
timestamp 1644511149
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_641
timestamp 1644511149
transform 1 0 60076 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_668
timestamp 1644511149
transform 1 0 62560 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_673
timestamp 1644511149
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_685
timestamp 1644511149
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_697
timestamp 1644511149
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_709
timestamp 1644511149
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1644511149
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1644511149
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_729
timestamp 1644511149
transform 1 0 68172 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_295
timestamp 1644511149
transform 1 0 28244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_355
timestamp 1644511149
transform 1 0 33764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_541
timestamp 1644511149
transform 1 0 50876 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_564
timestamp 1644511149
transform 1 0 52992 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_576
timestamp 1644511149
transform 1 0 54096 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_601
timestamp 1644511149
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_613
timestamp 1644511149
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_625
timestamp 1644511149
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1644511149
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1644511149
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_645
timestamp 1644511149
transform 1 0 60444 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_656
timestamp 1644511149
transform 1 0 61456 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_668
timestamp 1644511149
transform 1 0 62560 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_680
timestamp 1644511149
transform 1 0 63664 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_692
timestamp 1644511149
transform 1 0 64768 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_701
timestamp 1644511149
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_713
timestamp 1644511149
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_725
timestamp 1644511149
transform 1 0 67804 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_308
timestamp 1644511149
transform 1 0 29440 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_320
timestamp 1644511149
transform 1 0 30544 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_402
timestamp 1644511149
transform 1 0 38088 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_415
timestamp 1644511149
transform 1 0 39284 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_427
timestamp 1644511149
transform 1 0 40388 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_439
timestamp 1644511149
transform 1 0 41492 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_537
timestamp 1644511149
transform 1 0 50508 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_543
timestamp 1644511149
transform 1 0 51060 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_550
timestamp 1644511149
transform 1 0 51704 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_558
timestamp 1644511149
transform 1 0 52440 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1644511149
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1644511149
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_629
timestamp 1644511149
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_641
timestamp 1644511149
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_653
timestamp 1644511149
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1644511149
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1644511149
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_673
timestamp 1644511149
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_685
timestamp 1644511149
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_697
timestamp 1644511149
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_709
timestamp 1644511149
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1644511149
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1644511149
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_729
timestamp 1644511149
transform 1 0 68172 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1644511149
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_203
timestamp 1644511149
transform 1 0 19780 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_207
timestamp 1644511149
transform 1 0 20148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_219
timestamp 1644511149
transform 1 0 21252 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_231
timestamp 1644511149
transform 1 0 22356 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_243
timestamp 1644511149
transform 1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_286
timestamp 1644511149
transform 1 0 27416 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_294
timestamp 1644511149
transform 1 0 28152 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_298
timestamp 1644511149
transform 1 0 28520 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1644511149
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1644511149
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_544
timestamp 1644511149
transform 1 0 51152 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_625
timestamp 1644511149
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1644511149
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1644511149
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_645
timestamp 1644511149
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_657
timestamp 1644511149
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_669
timestamp 1644511149
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_681
timestamp 1644511149
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1644511149
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1644511149
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_701
timestamp 1644511149
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_713
timestamp 1644511149
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_725
timestamp 1644511149
transform 1 0 67804 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_266
timestamp 1644511149
transform 1 0 25576 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_288
timestamp 1644511149
transform 1 0 27600 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_313
timestamp 1644511149
transform 1 0 29900 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_325
timestamp 1644511149
transform 1 0 31004 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1644511149
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_547
timestamp 1644511149
transform 1 0 51428 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_629
timestamp 1644511149
transform 1 0 58972 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_637
timestamp 1644511149
transform 1 0 59708 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_643
timestamp 1644511149
transform 1 0 60260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_655
timestamp 1644511149
transform 1 0 61364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_667
timestamp 1644511149
transform 1 0 62468 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1644511149
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_673
timestamp 1644511149
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_685
timestamp 1644511149
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_697
timestamp 1644511149
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_709
timestamp 1644511149
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1644511149
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1644511149
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_729
timestamp 1644511149
transform 1 0 68172 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_68
timestamp 1644511149
transform 1 0 7360 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_72
timestamp 1644511149
transform 1 0 7728 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_76
timestamp 1644511149
transform 1 0 8096 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_203
timestamp 1644511149
transform 1 0 19780 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_215
timestamp 1644511149
transform 1 0 20884 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_227
timestamp 1644511149
transform 1 0 21988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_239
timestamp 1644511149
transform 1 0 23092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_296
timestamp 1644511149
transform 1 0 28336 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_341
timestamp 1644511149
transform 1 0 32476 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_353
timestamp 1644511149
transform 1 0 33580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1644511149
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_625
timestamp 1644511149
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_640
timestamp 1644511149
transform 1 0 59984 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_666
timestamp 1644511149
transform 1 0 62376 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_678
timestamp 1644511149
transform 1 0 63480 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_690
timestamp 1644511149
transform 1 0 64584 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_698
timestamp 1644511149
transform 1 0 65320 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_701
timestamp 1644511149
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_713
timestamp 1644511149
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_725
timestamp 1644511149
transform 1 0 67804 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_60
timestamp 1644511149
transform 1 0 6624 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_72
timestamp 1644511149
transform 1 0 7728 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_84
timestamp 1644511149
transform 1 0 8832 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_96
timestamp 1644511149
transform 1 0 9936 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1644511149
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_401
timestamp 1644511149
transform 1 0 37996 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_412
timestamp 1644511149
transform 1 0 39008 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_424
timestamp 1644511149
transform 1 0 40112 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_436
timestamp 1644511149
transform 1 0 41216 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_629
timestamp 1644511149
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_641
timestamp 1644511149
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_653
timestamp 1644511149
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1644511149
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1644511149
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_673
timestamp 1644511149
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_685
timestamp 1644511149
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_697
timestamp 1644511149
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_709
timestamp 1644511149
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1644511149
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1644511149
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_729
timestamp 1644511149
transform 1 0 68172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_50
timestamp 1644511149
transform 1 0 5704 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_62
timestamp 1644511149
transform 1 0 6808 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_74
timestamp 1644511149
transform 1 0 7912 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1644511149
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_480
timestamp 1644511149
transform 1 0 45264 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_492
timestamp 1644511149
transform 1 0 46368 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_504
timestamp 1644511149
transform 1 0 47472 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_516
timestamp 1644511149
transform 1 0 48576 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_528
timestamp 1644511149
transform 1 0 49680 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_625
timestamp 1644511149
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1644511149
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1644511149
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_645
timestamp 1644511149
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_657
timestamp 1644511149
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_669
timestamp 1644511149
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_681
timestamp 1644511149
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1644511149
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1644511149
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_701
timestamp 1644511149
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_713
timestamp 1644511149
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_725
timestamp 1644511149
transform 1 0 67804 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_468
timestamp 1644511149
transform 1 0 44160 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_493
timestamp 1644511149
transform 1 0 46460 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_501
timestamp 1644511149
transform 1 0 47196 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_629
timestamp 1644511149
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_641
timestamp 1644511149
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_653
timestamp 1644511149
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1644511149
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1644511149
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_673
timestamp 1644511149
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_685
timestamp 1644511149
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_697
timestamp 1644511149
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_709
timestamp 1644511149
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 1644511149
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 1644511149
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_729
timestamp 1644511149
transform 1 0 68172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_448
timestamp 1644511149
transform 1 0 42320 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_460
timestamp 1644511149
transform 1 0 43424 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_472
timestamp 1644511149
transform 1 0 44528 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_513
timestamp 1644511149
transform 1 0 48300 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_524
timestamp 1644511149
transform 1 0 49312 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_600
timestamp 1644511149
transform 1 0 56304 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_612
timestamp 1644511149
transform 1 0 57408 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_624
timestamp 1644511149
transform 1 0 58512 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_636
timestamp 1644511149
transform 1 0 59616 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_645
timestamp 1644511149
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_657
timestamp 1644511149
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_669
timestamp 1644511149
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_681
timestamp 1644511149
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1644511149
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1644511149
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_701
timestamp 1644511149
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_713
timestamp 1644511149
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_725
timestamp 1644511149
transform 1 0 67804 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_264
timestamp 1644511149
transform 1 0 25392 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_444
timestamp 1644511149
transform 1 0 41952 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_470
timestamp 1644511149
transform 1 0 44344 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_482
timestamp 1644511149
transform 1 0 45448 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_494
timestamp 1644511149
transform 1 0 46552 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_502
timestamp 1644511149
transform 1 0 47288 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_521
timestamp 1644511149
transform 1 0 49036 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_543
timestamp 1644511149
transform 1 0 51060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_555
timestamp 1644511149
transform 1 0 52164 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_612
timestamp 1644511149
transform 1 0 57408 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_629
timestamp 1644511149
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_641
timestamp 1644511149
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_653
timestamp 1644511149
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1644511149
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1644511149
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_673
timestamp 1644511149
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_685
timestamp 1644511149
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_697
timestamp 1644511149
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_709
timestamp 1644511149
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 1644511149
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1644511149
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_729
timestamp 1644511149
transform 1 0 68172 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_257
timestamp 1644511149
transform 1 0 24748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_279
timestamp 1644511149
transform 1 0 26772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_291
timestamp 1644511149
transform 1 0 27876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_303
timestamp 1644511149
transform 1 0 28980 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_378
timestamp 1644511149
transform 1 0 35880 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_382
timestamp 1644511149
transform 1 0 36248 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_392
timestamp 1644511149
transform 1 0 37168 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_404
timestamp 1644511149
transform 1 0 38272 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_416
timestamp 1644511149
transform 1 0 39376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_513
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_521
timestamp 1644511149
transform 1 0 49036 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_526
timestamp 1644511149
transform 1 0 49496 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_598
timestamp 1644511149
transform 1 0 56120 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_610
timestamp 1644511149
transform 1 0 57224 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_622
timestamp 1644511149
transform 1 0 58328 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_634
timestamp 1644511149
transform 1 0 59432 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_642
timestamp 1644511149
transform 1 0 60168 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_645
timestamp 1644511149
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_657
timestamp 1644511149
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_669
timestamp 1644511149
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_681
timestamp 1644511149
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1644511149
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1644511149
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_701
timestamp 1644511149
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_713
timestamp 1644511149
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_725
timestamp 1644511149
transform 1 0 67804 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_257
timestamp 1644511149
transform 1 0 24748 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_381
timestamp 1644511149
transform 1 0 36156 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1644511149
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_402
timestamp 1644511149
transform 1 0 38088 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_414
timestamp 1644511149
transform 1 0 39192 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_426
timestamp 1644511149
transform 1 0 40296 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_438
timestamp 1644511149
transform 1 0 41400 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_446
timestamp 1644511149
transform 1 0 42136 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_517
timestamp 1644511149
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_529
timestamp 1644511149
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_541
timestamp 1644511149
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1644511149
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_629
timestamp 1644511149
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_641
timestamp 1644511149
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_653
timestamp 1644511149
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1644511149
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1644511149
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_673
timestamp 1644511149
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_685
timestamp 1644511149
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_697
timestamp 1644511149
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_709
timestamp 1644511149
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1644511149
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1644511149
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_729
timestamp 1644511149
transform 1 0 68172 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_60
timestamp 1644511149
transform 1 0 6624 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_72
timestamp 1644511149
transform 1 0 7728 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_513
timestamp 1644511149
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_625
timestamp 1644511149
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1644511149
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1644511149
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_645
timestamp 1644511149
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_657
timestamp 1644511149
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_669
timestamp 1644511149
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_681
timestamp 1644511149
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1644511149
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1644511149
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_701
timestamp 1644511149
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_713
timestamp 1644511149
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_725
timestamp 1644511149
transform 1 0 67804 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_78
timestamp 1644511149
transform 1 0 8280 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_90
timestamp 1644511149
transform 1 0 9384 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_102
timestamp 1644511149
transform 1 0 10488 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1644511149
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_347
timestamp 1644511149
transform 1 0 33028 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_355
timestamp 1644511149
transform 1 0 33764 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_365
timestamp 1644511149
transform 1 0 34684 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_381
timestamp 1644511149
transform 1 0 36156 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_389
timestamp 1644511149
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_469
timestamp 1644511149
transform 1 0 44252 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_475
timestamp 1644511149
transform 1 0 44804 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_500
timestamp 1644511149
transform 1 0 47104 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_529
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_541
timestamp 1644511149
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1644511149
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_629
timestamp 1644511149
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_641
timestamp 1644511149
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_653
timestamp 1644511149
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1644511149
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1644511149
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_673
timestamp 1644511149
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_685
timestamp 1644511149
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_697
timestamp 1644511149
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_709
timestamp 1644511149
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1644511149
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1644511149
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_729
timestamp 1644511149
transform 1 0 68172 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_58
timestamp 1644511149
transform 1 0 6440 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_70
timestamp 1644511149
transform 1 0 7544 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1644511149
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_144
timestamp 1644511149
transform 1 0 14352 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_156
timestamp 1644511149
transform 1 0 15456 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_168
timestamp 1644511149
transform 1 0 16560 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_180
timestamp 1644511149
transform 1 0 17664 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_348
timestamp 1644511149
transform 1 0 33120 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_358
timestamp 1644511149
transform 1 0 34040 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_381
timestamp 1644511149
transform 1 0 36156 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_404
timestamp 1644511149
transform 1 0 38272 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_416
timestamp 1644511149
transform 1 0 39376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_484
timestamp 1644511149
transform 1 0 45632 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_496
timestamp 1644511149
transform 1 0 46736 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_508
timestamp 1644511149
transform 1 0 47840 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_520
timestamp 1644511149
transform 1 0 48944 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_625
timestamp 1644511149
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1644511149
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1644511149
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_645
timestamp 1644511149
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_657
timestamp 1644511149
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_669
timestamp 1644511149
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_681
timestamp 1644511149
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1644511149
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1644511149
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_722
timestamp 1644511149
transform 1 0 67528 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_730
timestamp 1644511149
transform 1 0 68264 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_131
timestamp 1644511149
transform 1 0 13156 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_135
timestamp 1644511149
transform 1 0 13524 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_160
timestamp 1644511149
transform 1 0 15824 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_345
timestamp 1644511149
transform 1 0 32844 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_353
timestamp 1644511149
transform 1 0 33580 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_366
timestamp 1644511149
transform 1 0 34776 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_379
timestamp 1644511149
transform 1 0 35972 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1644511149
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_402
timestamp 1644511149
transform 1 0 38088 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_415
timestamp 1644511149
transform 1 0 39284 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_428
timestamp 1644511149
transform 1 0 40480 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_440
timestamp 1644511149
transform 1 0 41584 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_629
timestamp 1644511149
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_641
timestamp 1644511149
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_653
timestamp 1644511149
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1644511149
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1644511149
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_673
timestamp 1644511149
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_685
timestamp 1644511149
transform 1 0 64124 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_691
timestamp 1644511149
transform 1 0 64676 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_695
timestamp 1644511149
transform 1 0 65044 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_702
timestamp 1644511149
transform 1 0 65688 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_714
timestamp 1644511149
transform 1 0 66792 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_726
timestamp 1644511149
transform 1 0 67896 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_729
timestamp 1644511149
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_343
timestamp 1644511149
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_355
timestamp 1644511149
transform 1 0 33764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_371
timestamp 1644511149
transform 1 0 35236 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_376
timestamp 1644511149
transform 1 0 35696 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_388
timestamp 1644511149
transform 1 0 36800 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_415
timestamp 1644511149
transform 1 0 39284 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1644511149
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1644511149
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_545
timestamp 1644511149
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_557
timestamp 1644511149
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_569
timestamp 1644511149
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1644511149
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1644511149
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_601
timestamp 1644511149
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_613
timestamp 1644511149
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_625
timestamp 1644511149
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_637
timestamp 1644511149
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1644511149
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_645
timestamp 1644511149
transform 1 0 60444 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_654
timestamp 1644511149
transform 1 0 61272 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_679
timestamp 1644511149
transform 1 0 63572 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_691
timestamp 1644511149
transform 1 0 64676 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_699
timestamp 1644511149
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_701
timestamp 1644511149
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_713
timestamp 1644511149
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_725
timestamp 1644511149
transform 1 0 67804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_397
timestamp 1644511149
transform 1 0 37628 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_409
timestamp 1644511149
transform 1 0 38732 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_421
timestamp 1644511149
transform 1 0 39836 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_433
timestamp 1644511149
transform 1 0 40940 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_445
timestamp 1644511149
transform 1 0 42044 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_517
timestamp 1644511149
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_529
timestamp 1644511149
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_541
timestamp 1644511149
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1644511149
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1644511149
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_561
timestamp 1644511149
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_573
timestamp 1644511149
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_585
timestamp 1644511149
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_597
timestamp 1644511149
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1644511149
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1644511149
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_617
timestamp 1644511149
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_629
timestamp 1644511149
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_641
timestamp 1644511149
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_653
timestamp 1644511149
transform 1 0 61180 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_657
timestamp 1644511149
transform 1 0 61548 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_661
timestamp 1644511149
transform 1 0 61916 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_669
timestamp 1644511149
transform 1 0 62652 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_673
timestamp 1644511149
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_685
timestamp 1644511149
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_697
timestamp 1644511149
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_709
timestamp 1644511149
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_721
timestamp 1644511149
transform 1 0 67436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_727
timestamp 1644511149
transform 1 0 67988 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_729
timestamp 1644511149
transform 1 0 68172 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_348
timestamp 1644511149
transform 1 0 33120 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_360
timestamp 1644511149
transform 1 0 34224 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_501
timestamp 1644511149
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_513
timestamp 1644511149
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1644511149
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1644511149
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_533
timestamp 1644511149
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_545
timestamp 1644511149
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_557
timestamp 1644511149
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_569
timestamp 1644511149
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1644511149
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1644511149
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_589
timestamp 1644511149
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_601
timestamp 1644511149
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_613
timestamp 1644511149
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_625
timestamp 1644511149
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_637
timestamp 1644511149
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_643
timestamp 1644511149
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_645
timestamp 1644511149
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_657
timestamp 1644511149
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_669
timestamp 1644511149
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_681
timestamp 1644511149
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_693
timestamp 1644511149
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_699
timestamp 1644511149
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_704
timestamp 1644511149
transform 1 0 65872 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_716
timestamp 1644511149
transform 1 0 66976 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_728
timestamp 1644511149
transform 1 0 68080 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_732
timestamp 1644511149
transform 1 0 68448 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_99
timestamp 1644511149
transform 1 0 10212 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_103
timestamp 1644511149
transform 1 0 10580 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_345
timestamp 1644511149
transform 1 0 32844 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_367
timestamp 1644511149
transform 1 0 34868 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_379
timestamp 1644511149
transform 1 0 35972 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_517
timestamp 1644511149
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_529
timestamp 1644511149
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_541
timestamp 1644511149
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1644511149
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1644511149
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_561
timestamp 1644511149
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_573
timestamp 1644511149
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_585
timestamp 1644511149
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_597
timestamp 1644511149
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1644511149
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1644511149
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_617
timestamp 1644511149
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_629
timestamp 1644511149
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_641
timestamp 1644511149
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_653
timestamp 1644511149
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1644511149
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1644511149
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_673
timestamp 1644511149
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_685
timestamp 1644511149
transform 1 0 64124 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_694
timestamp 1644511149
transform 1 0 64952 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_719
timestamp 1644511149
transform 1 0 67252 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_727
timestamp 1644511149
transform 1 0 67988 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_729
timestamp 1644511149
transform 1 0 68172 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_93
timestamp 1644511149
transform 1 0 9660 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_115
timestamp 1644511149
transform 1 0 11684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_127
timestamp 1644511149
transform 1 0 12788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_350
timestamp 1644511149
transform 1 0 33304 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_362
timestamp 1644511149
transform 1 0 34408 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_501
timestamp 1644511149
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_513
timestamp 1644511149
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1644511149
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1644511149
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_533
timestamp 1644511149
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_545
timestamp 1644511149
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_557
timestamp 1644511149
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_569
timestamp 1644511149
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1644511149
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1644511149
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_589
timestamp 1644511149
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_601
timestamp 1644511149
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_613
timestamp 1644511149
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_625
timestamp 1644511149
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_637
timestamp 1644511149
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1644511149
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_645
timestamp 1644511149
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_657
timestamp 1644511149
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_669
timestamp 1644511149
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_681
timestamp 1644511149
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1644511149
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1644511149
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_701
timestamp 1644511149
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_713
timestamp 1644511149
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_725
timestamp 1644511149
transform 1 0 67804 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_98
timestamp 1644511149
transform 1 0 10120 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_110
timestamp 1644511149
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_505
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_517
timestamp 1644511149
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_529
timestamp 1644511149
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_541
timestamp 1644511149
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1644511149
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1644511149
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_561
timestamp 1644511149
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_573
timestamp 1644511149
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_585
timestamp 1644511149
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_597
timestamp 1644511149
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1644511149
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1644511149
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_617
timestamp 1644511149
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_629
timestamp 1644511149
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_641
timestamp 1644511149
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_653
timestamp 1644511149
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_665
timestamp 1644511149
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_671
timestamp 1644511149
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_673
timestamp 1644511149
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_685
timestamp 1644511149
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_697
timestamp 1644511149
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_709
timestamp 1644511149
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_721
timestamp 1644511149
transform 1 0 67436 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_727
timestamp 1644511149
transform 1 0 67988 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_729
timestamp 1644511149
transform 1 0 68172 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_513
timestamp 1644511149
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1644511149
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1644511149
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_533
timestamp 1644511149
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_545
timestamp 1644511149
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_557
timestamp 1644511149
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_569
timestamp 1644511149
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1644511149
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1644511149
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_589
timestamp 1644511149
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_601
timestamp 1644511149
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_613
timestamp 1644511149
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_625
timestamp 1644511149
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_637
timestamp 1644511149
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1644511149
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_645
timestamp 1644511149
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_657
timestamp 1644511149
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_669
timestamp 1644511149
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_681
timestamp 1644511149
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1644511149
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1644511149
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_701
timestamp 1644511149
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_713
timestamp 1644511149
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_725
timestamp 1644511149
transform 1 0 67804 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1644511149
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1644511149
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_517
timestamp 1644511149
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_529
timestamp 1644511149
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_541
timestamp 1644511149
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1644511149
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1644511149
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_561
timestamp 1644511149
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_573
timestamp 1644511149
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_585
timestamp 1644511149
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_597
timestamp 1644511149
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1644511149
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1644511149
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_617
timestamp 1644511149
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_629
timestamp 1644511149
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_641
timestamp 1644511149
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_653
timestamp 1644511149
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1644511149
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_671
timestamp 1644511149
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_673
timestamp 1644511149
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_685
timestamp 1644511149
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_697
timestamp 1644511149
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_709
timestamp 1644511149
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_721
timestamp 1644511149
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_727
timestamp 1644511149
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_729
timestamp 1644511149
transform 1 0 68172 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_501
timestamp 1644511149
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_513
timestamp 1644511149
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1644511149
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1644511149
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_533
timestamp 1644511149
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_545
timestamp 1644511149
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_557
timestamp 1644511149
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_569
timestamp 1644511149
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1644511149
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1644511149
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_589
timestamp 1644511149
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_601
timestamp 1644511149
transform 1 0 56396 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_608
timestamp 1644511149
transform 1 0 57040 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_633
timestamp 1644511149
transform 1 0 59340 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_641
timestamp 1644511149
transform 1 0 60076 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_645
timestamp 1644511149
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_657
timestamp 1644511149
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_669
timestamp 1644511149
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_681
timestamp 1644511149
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1644511149
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1644511149
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_701
timestamp 1644511149
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_713
timestamp 1644511149
transform 1 0 66700 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_725
timestamp 1644511149
transform 1 0 67804 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1644511149
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1644511149
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_174
timestamp 1644511149
transform 1 0 17112 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_186
timestamp 1644511149
transform 1 0 18216 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_198
timestamp 1644511149
transform 1 0 19320 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_210
timestamp 1644511149
transform 1 0 20424 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1644511149
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_366
timestamp 1644511149
transform 1 0 34776 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_378
timestamp 1644511149
transform 1 0 35880 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_390
timestamp 1644511149
transform 1 0 36984 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_479
timestamp 1644511149
transform 1 0 45172 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_491
timestamp 1644511149
transform 1 0 46276 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1644511149
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_505
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_517
timestamp 1644511149
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_529
timestamp 1644511149
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_541
timestamp 1644511149
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1644511149
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1644511149
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_561
timestamp 1644511149
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_573
timestamp 1644511149
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_585
timestamp 1644511149
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_597
timestamp 1644511149
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1644511149
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1644511149
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_620
timestamp 1644511149
transform 1 0 58144 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_632
timestamp 1644511149
transform 1 0 59248 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_644
timestamp 1644511149
transform 1 0 60352 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_656
timestamp 1644511149
transform 1 0 61456 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_668
timestamp 1644511149
transform 1 0 62560 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_673
timestamp 1644511149
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_685
timestamp 1644511149
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_697
timestamp 1644511149
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_709
timestamp 1644511149
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_721
timestamp 1644511149
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_727
timestamp 1644511149
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_729
timestamp 1644511149
transform 1 0 68172 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_169
timestamp 1644511149
transform 1 0 16652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_191
timestamp 1644511149
transform 1 0 18676 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_386
timestamp 1644511149
transform 1 0 36616 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_398
timestamp 1644511149
transform 1 0 37720 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_410
timestamp 1644511149
transform 1 0 38824 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_418
timestamp 1644511149
transform 1 0 39560 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_498
timestamp 1644511149
transform 1 0 46920 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_510
timestamp 1644511149
transform 1 0 48024 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_522
timestamp 1644511149
transform 1 0 49128 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_530
timestamp 1644511149
transform 1 0 49864 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_533
timestamp 1644511149
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_545
timestamp 1644511149
transform 1 0 51244 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_551
timestamp 1644511149
transform 1 0 51796 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_576
timestamp 1644511149
transform 1 0 54096 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_589
timestamp 1644511149
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_601
timestamp 1644511149
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_613
timestamp 1644511149
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_625
timestamp 1644511149
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_637
timestamp 1644511149
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_643
timestamp 1644511149
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_648
timestamp 1644511149
transform 1 0 60720 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_660
timestamp 1644511149
transform 1 0 61824 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_672
timestamp 1644511149
transform 1 0 62928 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_684
timestamp 1644511149
transform 1 0 64032 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_696
timestamp 1644511149
transform 1 0 65136 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_701
timestamp 1644511149
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_713
timestamp 1644511149
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_725
timestamp 1644511149
transform 1 0 67804 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_174
timestamp 1644511149
transform 1 0 17112 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_186
timestamp 1644511149
transform 1 0 18216 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_198
timestamp 1644511149
transform 1 0 19320 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_210
timestamp 1644511149
transform 1 0 20424 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_222
timestamp 1644511149
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_360
timestamp 1644511149
transform 1 0 34224 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_372
timestamp 1644511149
transform 1 0 35328 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_384
timestamp 1644511149
transform 1 0 36432 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_477
timestamp 1644511149
transform 1 0 44988 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_481
timestamp 1644511149
transform 1 0 45356 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_493
timestamp 1644511149
transform 1 0 46460 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_501
timestamp 1644511149
transform 1 0 47196 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_505
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_517
timestamp 1644511149
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_529
timestamp 1644511149
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_541
timestamp 1644511149
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1644511149
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1644511149
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_564
timestamp 1644511149
transform 1 0 52992 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_576
timestamp 1644511149
transform 1 0 54096 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_588
timestamp 1644511149
transform 1 0 55200 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_600
timestamp 1644511149
transform 1 0 56304 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_612
timestamp 1644511149
transform 1 0 57408 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_617
timestamp 1644511149
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_629
timestamp 1644511149
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_641
timestamp 1644511149
transform 1 0 60076 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_664
timestamp 1644511149
transform 1 0 62192 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_673
timestamp 1644511149
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_685
timestamp 1644511149
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_697
timestamp 1644511149
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_709
timestamp 1644511149
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_721
timestamp 1644511149
transform 1 0 67436 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_727
timestamp 1644511149
transform 1 0 67988 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_729
timestamp 1644511149
transform 1 0 68172 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_489
timestamp 1644511149
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_501
timestamp 1644511149
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_513
timestamp 1644511149
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1644511149
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1644511149
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_533
timestamp 1644511149
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_545
timestamp 1644511149
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_557
timestamp 1644511149
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_569
timestamp 1644511149
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1644511149
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1644511149
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_589
timestamp 1644511149
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_601
timestamp 1644511149
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_613
timestamp 1644511149
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_625
timestamp 1644511149
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1644511149
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1644511149
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_648
timestamp 1644511149
transform 1 0 60720 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_660
timestamp 1644511149
transform 1 0 61824 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_672
timestamp 1644511149
transform 1 0 62928 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_684
timestamp 1644511149
transform 1 0 64032 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_696
timestamp 1644511149
transform 1 0 65136 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_701
timestamp 1644511149
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_713
timestamp 1644511149
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_725
timestamp 1644511149
transform 1 0 67804 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_485
timestamp 1644511149
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1644511149
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_505
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_517
timestamp 1644511149
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_529
timestamp 1644511149
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_541
timestamp 1644511149
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1644511149
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1644511149
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_561
timestamp 1644511149
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_573
timestamp 1644511149
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_585
timestamp 1644511149
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_597
timestamp 1644511149
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1644511149
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1644511149
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_617
timestamp 1644511149
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_629
timestamp 1644511149
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_641
timestamp 1644511149
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_653
timestamp 1644511149
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1644511149
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1644511149
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_673
timestamp 1644511149
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_685
timestamp 1644511149
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_697
timestamp 1644511149
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_709
timestamp 1644511149
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_721
timestamp 1644511149
transform 1 0 67436 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_727
timestamp 1644511149
transform 1 0 67988 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_729
timestamp 1644511149
transform 1 0 68172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_457
timestamp 1644511149
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1644511149
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_477
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_489
timestamp 1644511149
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_501
timestamp 1644511149
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_513
timestamp 1644511149
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1644511149
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1644511149
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_533
timestamp 1644511149
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_545
timestamp 1644511149
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_557
timestamp 1644511149
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_569
timestamp 1644511149
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1644511149
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1644511149
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_589
timestamp 1644511149
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_601
timestamp 1644511149
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_613
timestamp 1644511149
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_625
timestamp 1644511149
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1644511149
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1644511149
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_645
timestamp 1644511149
transform 1 0 60444 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_649
timestamp 1644511149
transform 1 0 60812 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_661
timestamp 1644511149
transform 1 0 61916 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_673
timestamp 1644511149
transform 1 0 63020 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_685
timestamp 1644511149
transform 1 0 64124 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_697
timestamp 1644511149
transform 1 0 65228 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_701
timestamp 1644511149
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_713
timestamp 1644511149
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_725
timestamp 1644511149
transform 1 0 67804 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1644511149
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1644511149
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1644511149
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_461
timestamp 1644511149
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_473
timestamp 1644511149
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_485
timestamp 1644511149
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1644511149
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_505
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_517
timestamp 1644511149
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_529
timestamp 1644511149
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_541
timestamp 1644511149
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1644511149
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1644511149
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_561
timestamp 1644511149
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_573
timestamp 1644511149
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_585
timestamp 1644511149
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_597
timestamp 1644511149
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1644511149
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1644511149
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_617
timestamp 1644511149
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_629
timestamp 1644511149
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_641
timestamp 1644511149
transform 1 0 60076 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_668
timestamp 1644511149
transform 1 0 62560 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_673
timestamp 1644511149
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_685
timestamp 1644511149
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_697
timestamp 1644511149
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_709
timestamp 1644511149
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_721
timestamp 1644511149
transform 1 0 67436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_727
timestamp 1644511149
transform 1 0 67988 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_729
timestamp 1644511149
transform 1 0 68172 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_221
timestamp 1644511149
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_233
timestamp 1644511149
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_289
timestamp 1644511149
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1644511149
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1644511149
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_440
timestamp 1644511149
transform 1 0 41584 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_465
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_473
timestamp 1644511149
transform 1 0 44620 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_489
timestamp 1644511149
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_501
timestamp 1644511149
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_513
timestamp 1644511149
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1644511149
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1644511149
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_533
timestamp 1644511149
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_545
timestamp 1644511149
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_557
timestamp 1644511149
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_569
timestamp 1644511149
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1644511149
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1644511149
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_589
timestamp 1644511149
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_601
timestamp 1644511149
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_613
timestamp 1644511149
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_625
timestamp 1644511149
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1644511149
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1644511149
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_645
timestamp 1644511149
transform 1 0 60444 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_654
timestamp 1644511149
transform 1 0 61272 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_666
timestamp 1644511149
transform 1 0 62376 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_678
timestamp 1644511149
transform 1 0 63480 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_690
timestamp 1644511149
transform 1 0 64584 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_698
timestamp 1644511149
transform 1 0 65320 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_701
timestamp 1644511149
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_713
timestamp 1644511149
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_725
timestamp 1644511149
transform 1 0 67804 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1644511149
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1644511149
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_205
timestamp 1644511149
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1644511149
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1644511149
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1644511149
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_405
timestamp 1644511149
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_417
timestamp 1644511149
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_429
timestamp 1644511149
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1644511149
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_452
timestamp 1644511149
transform 1 0 42688 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_464
timestamp 1644511149
transform 1 0 43792 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_476
timestamp 1644511149
transform 1 0 44896 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_488
timestamp 1644511149
transform 1 0 46000 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_517
timestamp 1644511149
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_529
timestamp 1644511149
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_541
timestamp 1644511149
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1644511149
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1644511149
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_561
timestamp 1644511149
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_573
timestamp 1644511149
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_585
timestamp 1644511149
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_597
timestamp 1644511149
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1644511149
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1644511149
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_617
timestamp 1644511149
transform 1 0 57868 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_621
timestamp 1644511149
transform 1 0 58236 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_633
timestamp 1644511149
transform 1 0 59340 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_645
timestamp 1644511149
transform 1 0 60444 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_657
timestamp 1644511149
transform 1 0 61548 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_661
timestamp 1644511149
transform 1 0 61916 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_669
timestamp 1644511149
transform 1 0 62652 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_673
timestamp 1644511149
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_685
timestamp 1644511149
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_697
timestamp 1644511149
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_709
timestamp 1644511149
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_721
timestamp 1644511149
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_727
timestamp 1644511149
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_729
timestamp 1644511149
transform 1 0 68172 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1644511149
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1644511149
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1644511149
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_121
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1644511149
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_177
timestamp 1644511149
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1644511149
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_209
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_221
timestamp 1644511149
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_233
timestamp 1644511149
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1644511149
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1644511149
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_289
timestamp 1644511149
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1644511149
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_333
timestamp 1644511149
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_345
timestamp 1644511149
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1644511149
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1644511149
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1644511149
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1644511149
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_433
timestamp 1644511149
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_445
timestamp 1644511149
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_457
timestamp 1644511149
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1644511149
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1644511149
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_489
timestamp 1644511149
transform 1 0 46092 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_512
timestamp 1644511149
transform 1 0 48208 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_524
timestamp 1644511149
transform 1 0 49312 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_533
timestamp 1644511149
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_545
timestamp 1644511149
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_557
timestamp 1644511149
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_569
timestamp 1644511149
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1644511149
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1644511149
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_589
timestamp 1644511149
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_601
timestamp 1644511149
transform 1 0 56396 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_609
timestamp 1644511149
transform 1 0 57132 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_613
timestamp 1644511149
transform 1 0 57500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_638
timestamp 1644511149
transform 1 0 59800 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_645
timestamp 1644511149
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_657
timestamp 1644511149
transform 1 0 61548 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_682
timestamp 1644511149
transform 1 0 63848 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_694
timestamp 1644511149
transform 1 0 64952 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_701
timestamp 1644511149
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_713
timestamp 1644511149
transform 1 0 66700 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_725
timestamp 1644511149
transform 1 0 67804 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1644511149
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1644511149
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_39
timestamp 1644511149
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1644511149
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1644511149
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1644511149
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1644511149
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_93
timestamp 1644511149
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1644511149
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1644511149
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_113
timestamp 1644511149
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_125
timestamp 1644511149
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_137
timestamp 1644511149
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_149
timestamp 1644511149
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1644511149
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1644511149
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_169
timestamp 1644511149
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_181
timestamp 1644511149
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_193
timestamp 1644511149
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_205
timestamp 1644511149
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1644511149
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1644511149
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_228
timestamp 1644511149
transform 1 0 22080 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_240
timestamp 1644511149
transform 1 0 23184 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_252
timestamp 1644511149
transform 1 0 24288 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_264
timestamp 1644511149
transform 1 0 25392 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_276
timestamp 1644511149
transform 1 0 26496 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_281
timestamp 1644511149
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_293
timestamp 1644511149
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_305
timestamp 1644511149
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_317
timestamp 1644511149
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1644511149
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1644511149
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_337
timestamp 1644511149
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_349
timestamp 1644511149
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_361
timestamp 1644511149
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_373
timestamp 1644511149
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1644511149
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1644511149
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_393
timestamp 1644511149
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_405
timestamp 1644511149
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_417
timestamp 1644511149
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_429
timestamp 1644511149
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1644511149
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1644511149
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_449
timestamp 1644511149
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_461
timestamp 1644511149
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_473
timestamp 1644511149
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_485
timestamp 1644511149
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_500
timestamp 1644511149
transform 1 0 47104 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_526
timestamp 1644511149
transform 1 0 49496 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_538
timestamp 1644511149
transform 1 0 50600 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_550
timestamp 1644511149
transform 1 0 51704 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_558
timestamp 1644511149
transform 1 0 52440 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_561
timestamp 1644511149
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_573
timestamp 1644511149
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_585
timestamp 1644511149
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_597
timestamp 1644511149
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1644511149
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1644511149
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_617
timestamp 1644511149
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_629
timestamp 1644511149
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_641
timestamp 1644511149
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_653
timestamp 1644511149
transform 1 0 61180 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_83_664
timestamp 1644511149
transform 1 0 62192 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_673
timestamp 1644511149
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_685
timestamp 1644511149
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_697
timestamp 1644511149
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_709
timestamp 1644511149
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_721
timestamp 1644511149
transform 1 0 67436 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_727
timestamp 1644511149
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_729
timestamp 1644511149
transform 1 0 68172 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1644511149
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1644511149
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1644511149
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1644511149
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1644511149
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1644511149
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1644511149
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_97
timestamp 1644511149
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_109
timestamp 1644511149
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_121
timestamp 1644511149
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1644511149
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1644511149
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_141
timestamp 1644511149
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_153
timestamp 1644511149
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_165
timestamp 1644511149
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_177
timestamp 1644511149
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1644511149
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1644511149
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_197
timestamp 1644511149
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_209
timestamp 1644511149
transform 1 0 20332 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_213
timestamp 1644511149
transform 1 0 20700 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_235
timestamp 1644511149
transform 1 0 22724 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_247
timestamp 1644511149
transform 1 0 23828 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1644511149
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_253
timestamp 1644511149
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_265
timestamp 1644511149
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_277
timestamp 1644511149
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_289
timestamp 1644511149
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1644511149
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1644511149
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_309
timestamp 1644511149
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_321
timestamp 1644511149
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_333
timestamp 1644511149
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_345
timestamp 1644511149
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1644511149
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1644511149
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_365
timestamp 1644511149
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_377
timestamp 1644511149
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_389
timestamp 1644511149
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_401
timestamp 1644511149
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1644511149
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1644511149
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_421
timestamp 1644511149
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_433
timestamp 1644511149
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_445
timestamp 1644511149
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_457
timestamp 1644511149
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1644511149
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1644511149
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_477
timestamp 1644511149
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_489
timestamp 1644511149
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_501
timestamp 1644511149
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_513
timestamp 1644511149
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1644511149
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1644511149
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_533
timestamp 1644511149
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_545
timestamp 1644511149
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_557
timestamp 1644511149
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_569
timestamp 1644511149
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1644511149
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1644511149
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_589
timestamp 1644511149
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_601
timestamp 1644511149
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_613
timestamp 1644511149
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_625
timestamp 1644511149
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1644511149
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1644511149
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_645
timestamp 1644511149
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_657
timestamp 1644511149
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_669
timestamp 1644511149
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_681
timestamp 1644511149
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1644511149
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1644511149
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_701
timestamp 1644511149
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_713
timestamp 1644511149
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_725
timestamp 1644511149
transform 1 0 67804 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1644511149
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1644511149
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1644511149
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1644511149
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1644511149
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1644511149
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1644511149
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_93
timestamp 1644511149
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1644511149
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1644511149
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_113
timestamp 1644511149
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_125
timestamp 1644511149
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_137
timestamp 1644511149
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_149
timestamp 1644511149
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1644511149
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1644511149
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_169
timestamp 1644511149
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_181
timestamp 1644511149
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_193
timestamp 1644511149
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_205
timestamp 1644511149
transform 1 0 19964 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_213
timestamp 1644511149
transform 1 0 20700 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1644511149
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1644511149
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_225
timestamp 1644511149
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_237
timestamp 1644511149
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_249
timestamp 1644511149
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_261
timestamp 1644511149
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1644511149
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1644511149
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_281
timestamp 1644511149
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_293
timestamp 1644511149
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_305
timestamp 1644511149
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_317
timestamp 1644511149
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1644511149
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1644511149
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_337
timestamp 1644511149
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_349
timestamp 1644511149
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_361
timestamp 1644511149
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_373
timestamp 1644511149
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1644511149
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1644511149
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_393
timestamp 1644511149
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_405
timestamp 1644511149
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_417
timestamp 1644511149
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_429
timestamp 1644511149
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1644511149
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1644511149
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_449
timestamp 1644511149
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_461
timestamp 1644511149
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_473
timestamp 1644511149
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_485
timestamp 1644511149
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1644511149
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1644511149
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_505
timestamp 1644511149
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_517
timestamp 1644511149
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_529
timestamp 1644511149
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_541
timestamp 1644511149
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1644511149
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1644511149
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_561
timestamp 1644511149
transform 1 0 52716 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_85_572
timestamp 1644511149
transform 1 0 53728 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_597
timestamp 1644511149
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1644511149
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1644511149
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_617
timestamp 1644511149
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_629
timestamp 1644511149
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_641
timestamp 1644511149
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_653
timestamp 1644511149
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1644511149
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1644511149
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_673
timestamp 1644511149
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_685
timestamp 1644511149
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_697
timestamp 1644511149
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_709
timestamp 1644511149
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_721
timestamp 1644511149
transform 1 0 67436 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_727
timestamp 1644511149
transform 1 0 67988 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_729
timestamp 1644511149
transform 1 0 68172 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1644511149
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1644511149
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_41
timestamp 1644511149
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_53
timestamp 1644511149
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_65
timestamp 1644511149
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1644511149
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1644511149
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_85
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_97
timestamp 1644511149
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_109
timestamp 1644511149
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_121
timestamp 1644511149
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1644511149
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1644511149
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_141
timestamp 1644511149
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_153
timestamp 1644511149
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_165
timestamp 1644511149
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_177
timestamp 1644511149
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1644511149
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1644511149
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_197
timestamp 1644511149
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_209
timestamp 1644511149
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_221
timestamp 1644511149
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_233
timestamp 1644511149
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1644511149
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1644511149
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_253
timestamp 1644511149
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_265
timestamp 1644511149
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_277
timestamp 1644511149
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_289
timestamp 1644511149
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1644511149
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1644511149
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_309
timestamp 1644511149
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_321
timestamp 1644511149
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_333
timestamp 1644511149
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_345
timestamp 1644511149
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1644511149
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1644511149
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_365
timestamp 1644511149
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_377
timestamp 1644511149
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_389
timestamp 1644511149
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_401
timestamp 1644511149
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1644511149
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1644511149
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_421
timestamp 1644511149
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_433
timestamp 1644511149
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_445
timestamp 1644511149
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_457
timestamp 1644511149
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1644511149
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1644511149
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_477
timestamp 1644511149
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_489
timestamp 1644511149
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_501
timestamp 1644511149
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_513
timestamp 1644511149
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1644511149
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1644511149
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_533
timestamp 1644511149
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_545
timestamp 1644511149
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_557
timestamp 1644511149
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_569
timestamp 1644511149
transform 1 0 53452 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_86_580
timestamp 1644511149
transform 1 0 54464 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_589
timestamp 1644511149
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_601
timestamp 1644511149
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_613
timestamp 1644511149
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_625
timestamp 1644511149
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1644511149
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1644511149
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_645
timestamp 1644511149
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_657
timestamp 1644511149
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_669
timestamp 1644511149
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_681
timestamp 1644511149
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1644511149
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1644511149
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_701
timestamp 1644511149
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_713
timestamp 1644511149
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_725
timestamp 1644511149
transform 1 0 67804 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1644511149
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1644511149
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1644511149
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1644511149
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1644511149
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1644511149
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1644511149
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1644511149
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1644511149
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_93
timestamp 1644511149
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1644511149
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1644511149
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_113
timestamp 1644511149
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_125
timestamp 1644511149
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_137
timestamp 1644511149
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_149
timestamp 1644511149
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1644511149
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1644511149
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_169
timestamp 1644511149
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_181
timestamp 1644511149
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_193
timestamp 1644511149
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_205
timestamp 1644511149
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1644511149
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1644511149
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_225
timestamp 1644511149
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_237
timestamp 1644511149
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_249
timestamp 1644511149
transform 1 0 24012 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_260
timestamp 1644511149
transform 1 0 25024 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_272
timestamp 1644511149
transform 1 0 26128 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_281
timestamp 1644511149
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_293
timestamp 1644511149
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_305
timestamp 1644511149
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_317
timestamp 1644511149
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1644511149
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1644511149
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_337
timestamp 1644511149
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_349
timestamp 1644511149
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_361
timestamp 1644511149
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_373
timestamp 1644511149
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1644511149
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1644511149
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_393
timestamp 1644511149
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_405
timestamp 1644511149
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_417
timestamp 1644511149
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_429
timestamp 1644511149
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1644511149
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1644511149
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_449
timestamp 1644511149
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_461
timestamp 1644511149
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_473
timestamp 1644511149
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_485
timestamp 1644511149
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1644511149
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1644511149
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_505
timestamp 1644511149
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_517
timestamp 1644511149
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_529
timestamp 1644511149
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_541
timestamp 1644511149
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1644511149
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1644511149
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_561
timestamp 1644511149
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_573
timestamp 1644511149
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_585
timestamp 1644511149
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_597
timestamp 1644511149
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1644511149
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1644511149
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_617
timestamp 1644511149
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_629
timestamp 1644511149
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_641
timestamp 1644511149
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_653
timestamp 1644511149
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1644511149
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1644511149
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_673
timestamp 1644511149
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_685
timestamp 1644511149
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_697
timestamp 1644511149
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_709
timestamp 1644511149
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_721
timestamp 1644511149
transform 1 0 67436 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_727
timestamp 1644511149
transform 1 0 67988 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_729
timestamp 1644511149
transform 1 0 68172 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1644511149
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1644511149
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1644511149
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_29
timestamp 1644511149
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_41
timestamp 1644511149
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_53
timestamp 1644511149
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_65
timestamp 1644511149
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1644511149
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1644511149
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_85
timestamp 1644511149
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_97
timestamp 1644511149
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_109
timestamp 1644511149
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_121
timestamp 1644511149
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1644511149
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1644511149
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_141
timestamp 1644511149
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_153
timestamp 1644511149
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_165
timestamp 1644511149
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_177
timestamp 1644511149
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1644511149
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1644511149
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_197
timestamp 1644511149
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_209
timestamp 1644511149
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_221
timestamp 1644511149
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_233
timestamp 1644511149
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1644511149
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1644511149
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_274
timestamp 1644511149
transform 1 0 26312 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_286
timestamp 1644511149
transform 1 0 27416 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_298
timestamp 1644511149
transform 1 0 28520 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_306
timestamp 1644511149
transform 1 0 29256 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_88_309
timestamp 1644511149
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_321
timestamp 1644511149
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_333
timestamp 1644511149
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_345
timestamp 1644511149
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1644511149
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1644511149
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_365
timestamp 1644511149
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_377
timestamp 1644511149
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_389
timestamp 1644511149
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_401
timestamp 1644511149
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1644511149
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1644511149
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_421
timestamp 1644511149
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_433
timestamp 1644511149
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_445
timestamp 1644511149
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_457
timestamp 1644511149
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1644511149
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1644511149
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_477
timestamp 1644511149
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_489
timestamp 1644511149
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_501
timestamp 1644511149
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_513
timestamp 1644511149
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1644511149
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1644511149
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_533
timestamp 1644511149
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_545
timestamp 1644511149
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_557
timestamp 1644511149
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_569
timestamp 1644511149
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1644511149
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1644511149
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_589
timestamp 1644511149
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_601
timestamp 1644511149
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_613
timestamp 1644511149
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_625
timestamp 1644511149
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1644511149
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1644511149
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_645
timestamp 1644511149
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_657
timestamp 1644511149
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_669
timestamp 1644511149
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_681
timestamp 1644511149
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_693
timestamp 1644511149
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_699
timestamp 1644511149
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_701
timestamp 1644511149
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_713
timestamp 1644511149
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_725
timestamp 1644511149
transform 1 0 67804 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1644511149
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1644511149
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1644511149
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_39
timestamp 1644511149
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1644511149
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1644511149
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1644511149
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1644511149
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1644511149
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_93
timestamp 1644511149
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1644511149
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1644511149
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_113
timestamp 1644511149
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_125
timestamp 1644511149
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_137
timestamp 1644511149
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_149
timestamp 1644511149
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1644511149
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1644511149
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_169
timestamp 1644511149
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_181
timestamp 1644511149
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_193
timestamp 1644511149
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_205
timestamp 1644511149
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1644511149
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1644511149
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_225
timestamp 1644511149
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_237
timestamp 1644511149
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_249
timestamp 1644511149
transform 1 0 24012 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_255
timestamp 1644511149
transform 1 0 24564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_267
timestamp 1644511149
transform 1 0 25668 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1644511149
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_281
timestamp 1644511149
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_293
timestamp 1644511149
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_305
timestamp 1644511149
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_317
timestamp 1644511149
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1644511149
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1644511149
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_337
timestamp 1644511149
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_349
timestamp 1644511149
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_361
timestamp 1644511149
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_373
timestamp 1644511149
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1644511149
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1644511149
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_393
timestamp 1644511149
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_405
timestamp 1644511149
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_417
timestamp 1644511149
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_429
timestamp 1644511149
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1644511149
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1644511149
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_449
timestamp 1644511149
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_461
timestamp 1644511149
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_473
timestamp 1644511149
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_485
timestamp 1644511149
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1644511149
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1644511149
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_505
timestamp 1644511149
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_517
timestamp 1644511149
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_529
timestamp 1644511149
transform 1 0 49772 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_537
timestamp 1644511149
transform 1 0 50508 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_542
timestamp 1644511149
transform 1 0 50968 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_554
timestamp 1644511149
transform 1 0 52072 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_561
timestamp 1644511149
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_573
timestamp 1644511149
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_585
timestamp 1644511149
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_597
timestamp 1644511149
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1644511149
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1644511149
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_617
timestamp 1644511149
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_629
timestamp 1644511149
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_641
timestamp 1644511149
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_653
timestamp 1644511149
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1644511149
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1644511149
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_673
timestamp 1644511149
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_685
timestamp 1644511149
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_697
timestamp 1644511149
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_709
timestamp 1644511149
transform 1 0 66332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_721
timestamp 1644511149
transform 1 0 67436 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_727
timestamp 1644511149
transform 1 0 67988 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_729
timestamp 1644511149
transform 1 0 68172 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1644511149
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1644511149
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1644511149
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1644511149
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1644511149
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1644511149
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1644511149
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1644511149
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1644511149
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_85
timestamp 1644511149
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_97
timestamp 1644511149
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_109
timestamp 1644511149
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_121
timestamp 1644511149
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1644511149
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1644511149
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_141
timestamp 1644511149
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_153
timestamp 1644511149
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_165
timestamp 1644511149
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_177
timestamp 1644511149
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1644511149
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1644511149
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_197
timestamp 1644511149
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_209
timestamp 1644511149
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_221
timestamp 1644511149
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_233
timestamp 1644511149
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1644511149
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1644511149
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_253
timestamp 1644511149
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_265
timestamp 1644511149
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_277
timestamp 1644511149
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_289
timestamp 1644511149
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1644511149
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1644511149
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_309
timestamp 1644511149
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_321
timestamp 1644511149
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_336
timestamp 1644511149
transform 1 0 32016 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_348
timestamp 1644511149
transform 1 0 33120 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_360
timestamp 1644511149
transform 1 0 34224 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_365
timestamp 1644511149
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_377
timestamp 1644511149
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_389
timestamp 1644511149
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_401
timestamp 1644511149
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1644511149
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1644511149
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_421
timestamp 1644511149
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_433
timestamp 1644511149
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_445
timestamp 1644511149
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_457
timestamp 1644511149
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1644511149
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1644511149
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_477
timestamp 1644511149
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_489
timestamp 1644511149
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_501
timestamp 1644511149
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_513
timestamp 1644511149
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1644511149
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1644511149
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_533
timestamp 1644511149
transform 1 0 50140 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_541
timestamp 1644511149
transform 1 0 50876 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_563
timestamp 1644511149
transform 1 0 52900 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_575
timestamp 1644511149
transform 1 0 54004 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1644511149
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_589
timestamp 1644511149
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_601
timestamp 1644511149
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_613
timestamp 1644511149
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_625
timestamp 1644511149
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1644511149
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1644511149
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_645
timestamp 1644511149
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_657
timestamp 1644511149
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_669
timestamp 1644511149
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_681
timestamp 1644511149
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1644511149
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1644511149
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_701
timestamp 1644511149
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_713
timestamp 1644511149
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_725
timestamp 1644511149
transform 1 0 67804 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1644511149
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_15
timestamp 1644511149
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_27
timestamp 1644511149
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_39
timestamp 1644511149
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1644511149
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1644511149
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1644511149
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1644511149
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1644511149
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_93
timestamp 1644511149
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1644511149
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1644511149
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_113
timestamp 1644511149
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_125
timestamp 1644511149
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_137
timestamp 1644511149
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_149
timestamp 1644511149
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1644511149
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1644511149
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_169
timestamp 1644511149
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_181
timestamp 1644511149
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_193
timestamp 1644511149
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_205
timestamp 1644511149
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1644511149
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1644511149
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_225
timestamp 1644511149
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_237
timestamp 1644511149
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_249
timestamp 1644511149
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_261
timestamp 1644511149
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1644511149
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1644511149
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_281
timestamp 1644511149
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_293
timestamp 1644511149
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_305
timestamp 1644511149
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_317
timestamp 1644511149
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_332
timestamp 1644511149
transform 1 0 31648 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_358
timestamp 1644511149
transform 1 0 34040 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_370
timestamp 1644511149
transform 1 0 35144 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_382
timestamp 1644511149
transform 1 0 36248 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_390
timestamp 1644511149
transform 1 0 36984 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_91_393
timestamp 1644511149
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_405
timestamp 1644511149
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_417
timestamp 1644511149
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_429
timestamp 1644511149
transform 1 0 40572 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_91_434
timestamp 1644511149
transform 1 0 41032 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_446
timestamp 1644511149
transform 1 0 42136 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_91_449
timestamp 1644511149
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_461
timestamp 1644511149
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_473
timestamp 1644511149
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_485
timestamp 1644511149
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1644511149
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1644511149
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_505
timestamp 1644511149
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_517
timestamp 1644511149
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_529
timestamp 1644511149
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_541
timestamp 1644511149
transform 1 0 50876 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_91_546
timestamp 1644511149
transform 1 0 51336 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_558
timestamp 1644511149
transform 1 0 52440 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_91_561
timestamp 1644511149
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_573
timestamp 1644511149
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_585
timestamp 1644511149
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_597
timestamp 1644511149
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1644511149
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1644511149
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_617
timestamp 1644511149
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_629
timestamp 1644511149
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_641
timestamp 1644511149
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_653
timestamp 1644511149
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1644511149
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1644511149
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_673
timestamp 1644511149
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_685
timestamp 1644511149
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_697
timestamp 1644511149
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_709
timestamp 1644511149
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_721
timestamp 1644511149
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_727
timestamp 1644511149
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_729
timestamp 1644511149
transform 1 0 68172 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1644511149
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1644511149
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1644511149
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1644511149
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1644511149
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1644511149
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1644511149
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1644511149
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1644511149
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_85
timestamp 1644511149
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_97
timestamp 1644511149
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_109
timestamp 1644511149
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_121
timestamp 1644511149
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1644511149
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1644511149
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_141
timestamp 1644511149
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_153
timestamp 1644511149
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_165
timestamp 1644511149
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_177
timestamp 1644511149
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1644511149
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1644511149
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_197
timestamp 1644511149
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_209
timestamp 1644511149
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_221
timestamp 1644511149
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_233
timestamp 1644511149
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1644511149
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1644511149
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_253
timestamp 1644511149
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_265
timestamp 1644511149
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_277
timestamp 1644511149
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_289
timestamp 1644511149
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1644511149
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1644511149
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_309
timestamp 1644511149
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_321
timestamp 1644511149
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_333
timestamp 1644511149
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_345
timestamp 1644511149
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1644511149
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1644511149
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_365
timestamp 1644511149
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_377
timestamp 1644511149
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_389
timestamp 1644511149
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_401
timestamp 1644511149
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1644511149
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1644511149
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_421
timestamp 1644511149
transform 1 0 39836 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_429
timestamp 1644511149
transform 1 0 40572 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_451
timestamp 1644511149
transform 1 0 42596 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_463
timestamp 1644511149
transform 1 0 43700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1644511149
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_477
timestamp 1644511149
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_489
timestamp 1644511149
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_501
timestamp 1644511149
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_513
timestamp 1644511149
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1644511149
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1644511149
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_533
timestamp 1644511149
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_545
timestamp 1644511149
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_557
timestamp 1644511149
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_569
timestamp 1644511149
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1644511149
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1644511149
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_589
timestamp 1644511149
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_601
timestamp 1644511149
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_613
timestamp 1644511149
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_625
timestamp 1644511149
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1644511149
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1644511149
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_645
timestamp 1644511149
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_657
timestamp 1644511149
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_669
timestamp 1644511149
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_681
timestamp 1644511149
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1644511149
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1644511149
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_701
timestamp 1644511149
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_713
timestamp 1644511149
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_725
timestamp 1644511149
transform 1 0 67804 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1644511149
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1644511149
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_27
timestamp 1644511149
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_39
timestamp 1644511149
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1644511149
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1644511149
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1644511149
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1644511149
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_81
timestamp 1644511149
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_93
timestamp 1644511149
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1644511149
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1644511149
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_113
timestamp 1644511149
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_125
timestamp 1644511149
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_137
timestamp 1644511149
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_149
timestamp 1644511149
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1644511149
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1644511149
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_169
timestamp 1644511149
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_181
timestamp 1644511149
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_193
timestamp 1644511149
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_205
timestamp 1644511149
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1644511149
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1644511149
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_225
timestamp 1644511149
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_237
timestamp 1644511149
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_249
timestamp 1644511149
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_261
timestamp 1644511149
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1644511149
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1644511149
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_281
timestamp 1644511149
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_293
timestamp 1644511149
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_305
timestamp 1644511149
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_317
timestamp 1644511149
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1644511149
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1644511149
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_337
timestamp 1644511149
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_349
timestamp 1644511149
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_361
timestamp 1644511149
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_373
timestamp 1644511149
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1644511149
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1644511149
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_393
timestamp 1644511149
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_405
timestamp 1644511149
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_417
timestamp 1644511149
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_429
timestamp 1644511149
transform 1 0 40572 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_434
timestamp 1644511149
transform 1 0 41032 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_446
timestamp 1644511149
transform 1 0 42136 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_449
timestamp 1644511149
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_461
timestamp 1644511149
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_473
timestamp 1644511149
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_485
timestamp 1644511149
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1644511149
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1644511149
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_505
timestamp 1644511149
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_517
timestamp 1644511149
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_529
timestamp 1644511149
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_541
timestamp 1644511149
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1644511149
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1644511149
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_561
timestamp 1644511149
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_573
timestamp 1644511149
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_585
timestamp 1644511149
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_597
timestamp 1644511149
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1644511149
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1644511149
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_617
timestamp 1644511149
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_629
timestamp 1644511149
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_641
timestamp 1644511149
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_653
timestamp 1644511149
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1644511149
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1644511149
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_673
timestamp 1644511149
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_685
timestamp 1644511149
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_697
timestamp 1644511149
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_709
timestamp 1644511149
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_721
timestamp 1644511149
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_727
timestamp 1644511149
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_729
timestamp 1644511149
transform 1 0 68172 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1644511149
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1644511149
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1644511149
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1644511149
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1644511149
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1644511149
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1644511149
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1644511149
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1644511149
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_85
timestamp 1644511149
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_97
timestamp 1644511149
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_109
timestamp 1644511149
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_121
timestamp 1644511149
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1644511149
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1644511149
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_141
timestamp 1644511149
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_153
timestamp 1644511149
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_165
timestamp 1644511149
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_177
timestamp 1644511149
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1644511149
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1644511149
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_197
timestamp 1644511149
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_209
timestamp 1644511149
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_221
timestamp 1644511149
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_233
timestamp 1644511149
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1644511149
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1644511149
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_253
timestamp 1644511149
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_265
timestamp 1644511149
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_277
timestamp 1644511149
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_289
timestamp 1644511149
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1644511149
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1644511149
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_309
timestamp 1644511149
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_321
timestamp 1644511149
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_333
timestamp 1644511149
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_345
timestamp 1644511149
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1644511149
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1644511149
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_365
timestamp 1644511149
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_377
timestamp 1644511149
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_389
timestamp 1644511149
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_401
timestamp 1644511149
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1644511149
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1644511149
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_421
timestamp 1644511149
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_433
timestamp 1644511149
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_445
timestamp 1644511149
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_457
timestamp 1644511149
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1644511149
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1644511149
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_477
timestamp 1644511149
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_489
timestamp 1644511149
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_501
timestamp 1644511149
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_513
timestamp 1644511149
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1644511149
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1644511149
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_533
timestamp 1644511149
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_545
timestamp 1644511149
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_557
timestamp 1644511149
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_569
timestamp 1644511149
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1644511149
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1644511149
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_589
timestamp 1644511149
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_601
timestamp 1644511149
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_613
timestamp 1644511149
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_625
timestamp 1644511149
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1644511149
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1644511149
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_645
timestamp 1644511149
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_657
timestamp 1644511149
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_669
timestamp 1644511149
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_681
timestamp 1644511149
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1644511149
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1644511149
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_701
timestamp 1644511149
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_713
timestamp 1644511149
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_725
timestamp 1644511149
transform 1 0 67804 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1644511149
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1644511149
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1644511149
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_39
timestamp 1644511149
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1644511149
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1644511149
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1644511149
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1644511149
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1644511149
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_93
timestamp 1644511149
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1644511149
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1644511149
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_113
timestamp 1644511149
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_125
timestamp 1644511149
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_137
timestamp 1644511149
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_149
timestamp 1644511149
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1644511149
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1644511149
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_169
timestamp 1644511149
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_181
timestamp 1644511149
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_193
timestamp 1644511149
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_205
timestamp 1644511149
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1644511149
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1644511149
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_225
timestamp 1644511149
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_237
timestamp 1644511149
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_249
timestamp 1644511149
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_261
timestamp 1644511149
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1644511149
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1644511149
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_281
timestamp 1644511149
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_293
timestamp 1644511149
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_305
timestamp 1644511149
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_317
timestamp 1644511149
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1644511149
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1644511149
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_337
timestamp 1644511149
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_349
timestamp 1644511149
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_361
timestamp 1644511149
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_373
timestamp 1644511149
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1644511149
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1644511149
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_393
timestamp 1644511149
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_405
timestamp 1644511149
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_417
timestamp 1644511149
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_429
timestamp 1644511149
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1644511149
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1644511149
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_449
timestamp 1644511149
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_461
timestamp 1644511149
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_473
timestamp 1644511149
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_485
timestamp 1644511149
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1644511149
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1644511149
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_505
timestamp 1644511149
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_517
timestamp 1644511149
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_529
timestamp 1644511149
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_541
timestamp 1644511149
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1644511149
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1644511149
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_561
timestamp 1644511149
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_573
timestamp 1644511149
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_585
timestamp 1644511149
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_597
timestamp 1644511149
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1644511149
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1644511149
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_617
timestamp 1644511149
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_629
timestamp 1644511149
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_641
timestamp 1644511149
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_653
timestamp 1644511149
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1644511149
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1644511149
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_673
timestamp 1644511149
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_685
timestamp 1644511149
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_697
timestamp 1644511149
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_709
timestamp 1644511149
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_721
timestamp 1644511149
transform 1 0 67436 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_727
timestamp 1644511149
transform 1 0 67988 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_729
timestamp 1644511149
transform 1 0 68172 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1644511149
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1644511149
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1644511149
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1644511149
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1644511149
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1644511149
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1644511149
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1644511149
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1644511149
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_85
timestamp 1644511149
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_97
timestamp 1644511149
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_109
timestamp 1644511149
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_121
timestamp 1644511149
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1644511149
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1644511149
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_141
timestamp 1644511149
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_153
timestamp 1644511149
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_165
timestamp 1644511149
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_177
timestamp 1644511149
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1644511149
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1644511149
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_197
timestamp 1644511149
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_209
timestamp 1644511149
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_221
timestamp 1644511149
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_233
timestamp 1644511149
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1644511149
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1644511149
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_253
timestamp 1644511149
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_265
timestamp 1644511149
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_277
timestamp 1644511149
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_289
timestamp 1644511149
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1644511149
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1644511149
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_309
timestamp 1644511149
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_321
timestamp 1644511149
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_333
timestamp 1644511149
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_345
timestamp 1644511149
transform 1 0 32844 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_351
timestamp 1644511149
transform 1 0 33396 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_355
timestamp 1644511149
transform 1 0 33764 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1644511149
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_368
timestamp 1644511149
transform 1 0 34960 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_380
timestamp 1644511149
transform 1 0 36064 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_392
timestamp 1644511149
transform 1 0 37168 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_404
timestamp 1644511149
transform 1 0 38272 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_416
timestamp 1644511149
transform 1 0 39376 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_421
timestamp 1644511149
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_433
timestamp 1644511149
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_445
timestamp 1644511149
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_457
timestamp 1644511149
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1644511149
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1644511149
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_477
timestamp 1644511149
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_489
timestamp 1644511149
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_501
timestamp 1644511149
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_513
timestamp 1644511149
transform 1 0 48300 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_519
timestamp 1644511149
transform 1 0 48852 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1644511149
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_533
timestamp 1644511149
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_545
timestamp 1644511149
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_557
timestamp 1644511149
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_569
timestamp 1644511149
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1644511149
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1644511149
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_589
timestamp 1644511149
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_601
timestamp 1644511149
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_613
timestamp 1644511149
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_625
timestamp 1644511149
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_637
timestamp 1644511149
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_643
timestamp 1644511149
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_645
timestamp 1644511149
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_657
timestamp 1644511149
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_669
timestamp 1644511149
transform 1 0 62652 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_96_696
timestamp 1644511149
transform 1 0 65136 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_701
timestamp 1644511149
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_713
timestamp 1644511149
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_725
timestamp 1644511149
transform 1 0 67804 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1644511149
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1644511149
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1644511149
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1644511149
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1644511149
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1644511149
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1644511149
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1644511149
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1644511149
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_93
timestamp 1644511149
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1644511149
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1644511149
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_113
timestamp 1644511149
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_125
timestamp 1644511149
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_137
timestamp 1644511149
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_149
timestamp 1644511149
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1644511149
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1644511149
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_169
timestamp 1644511149
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_181
timestamp 1644511149
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_193
timestamp 1644511149
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_205
timestamp 1644511149
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1644511149
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1644511149
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_225
timestamp 1644511149
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_237
timestamp 1644511149
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_249
timestamp 1644511149
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_261
timestamp 1644511149
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1644511149
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1644511149
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_281
timestamp 1644511149
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_293
timestamp 1644511149
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_305
timestamp 1644511149
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_317
timestamp 1644511149
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1644511149
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1644511149
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_337
timestamp 1644511149
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_349
timestamp 1644511149
transform 1 0 33212 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_373
timestamp 1644511149
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1644511149
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1644511149
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_393
timestamp 1644511149
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_405
timestamp 1644511149
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_417
timestamp 1644511149
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_429
timestamp 1644511149
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1644511149
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1644511149
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_449
timestamp 1644511149
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_461
timestamp 1644511149
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_473
timestamp 1644511149
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_485
timestamp 1644511149
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1644511149
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1644511149
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_505
timestamp 1644511149
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_538
timestamp 1644511149
transform 1 0 50600 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_550
timestamp 1644511149
transform 1 0 51704 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_558
timestamp 1644511149
transform 1 0 52440 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_561
timestamp 1644511149
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_573
timestamp 1644511149
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_585
timestamp 1644511149
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_597
timestamp 1644511149
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1644511149
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1644511149
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_617
timestamp 1644511149
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_629
timestamp 1644511149
transform 1 0 58972 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_641
timestamp 1644511149
transform 1 0 60076 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_653
timestamp 1644511149
transform 1 0 61180 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_665
timestamp 1644511149
transform 1 0 62284 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_671
timestamp 1644511149
transform 1 0 62836 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_97_673
timestamp 1644511149
transform 1 0 63020 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_679
timestamp 1644511149
transform 1 0 63572 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_683
timestamp 1644511149
transform 1 0 63940 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_691
timestamp 1644511149
transform 1 0 64676 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_715
timestamp 1644511149
transform 1 0 66884 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_727
timestamp 1644511149
transform 1 0 67988 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_729
timestamp 1644511149
transform 1 0 68172 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1644511149
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1644511149
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1644511149
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_29
timestamp 1644511149
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_41
timestamp 1644511149
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_53
timestamp 1644511149
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_65
timestamp 1644511149
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1644511149
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1644511149
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_85
timestamp 1644511149
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_97
timestamp 1644511149
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_109
timestamp 1644511149
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_121
timestamp 1644511149
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1644511149
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1644511149
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_141
timestamp 1644511149
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_153
timestamp 1644511149
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_165
timestamp 1644511149
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_177
timestamp 1644511149
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1644511149
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1644511149
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_197
timestamp 1644511149
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_209
timestamp 1644511149
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_221
timestamp 1644511149
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_233
timestamp 1644511149
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1644511149
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1644511149
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_253
timestamp 1644511149
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_265
timestamp 1644511149
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_277
timestamp 1644511149
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_289
timestamp 1644511149
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1644511149
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1644511149
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_309
timestamp 1644511149
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_321
timestamp 1644511149
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_333
timestamp 1644511149
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_345
timestamp 1644511149
transform 1 0 32844 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_349
timestamp 1644511149
transform 1 0 33212 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_356
timestamp 1644511149
transform 1 0 33856 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_365
timestamp 1644511149
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_377
timestamp 1644511149
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_389
timestamp 1644511149
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_401
timestamp 1644511149
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1644511149
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1644511149
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_421
timestamp 1644511149
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_433
timestamp 1644511149
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_445
timestamp 1644511149
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_457
timestamp 1644511149
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1644511149
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1644511149
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_477
timestamp 1644511149
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_489
timestamp 1644511149
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_501
timestamp 1644511149
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_98_513
timestamp 1644511149
transform 1 0 48300 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_518
timestamp 1644511149
transform 1 0 48760 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1644511149
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1644511149
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_533
timestamp 1644511149
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_545
timestamp 1644511149
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_557
timestamp 1644511149
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_569
timestamp 1644511149
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1644511149
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1644511149
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_589
timestamp 1644511149
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_601
timestamp 1644511149
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_613
timestamp 1644511149
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_625
timestamp 1644511149
transform 1 0 58604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_637
timestamp 1644511149
transform 1 0 59708 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_643
timestamp 1644511149
transform 1 0 60260 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_645
timestamp 1644511149
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_657
timestamp 1644511149
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_669
timestamp 1644511149
transform 1 0 62652 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_677
timestamp 1644511149
transform 1 0 63388 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_681
timestamp 1644511149
transform 1 0 63756 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_688
timestamp 1644511149
transform 1 0 64400 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_692
timestamp 1644511149
transform 1 0 64768 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_696
timestamp 1644511149
transform 1 0 65136 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_704
timestamp 1644511149
transform 1 0 65872 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_716
timestamp 1644511149
transform 1 0 66976 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_728
timestamp 1644511149
transform 1 0 68080 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_732
timestamp 1644511149
transform 1 0 68448 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1644511149
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1644511149
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_27
timestamp 1644511149
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_39
timestamp 1644511149
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1644511149
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1644511149
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1644511149
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1644511149
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1644511149
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_93
timestamp 1644511149
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1644511149
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1644511149
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_113
timestamp 1644511149
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_125
timestamp 1644511149
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_137
timestamp 1644511149
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_149
timestamp 1644511149
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1644511149
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1644511149
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_169
timestamp 1644511149
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_181
timestamp 1644511149
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_193
timestamp 1644511149
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_205
timestamp 1644511149
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1644511149
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1644511149
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_225
timestamp 1644511149
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_237
timestamp 1644511149
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_249
timestamp 1644511149
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_261
timestamp 1644511149
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1644511149
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1644511149
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_281
timestamp 1644511149
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_293
timestamp 1644511149
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_305
timestamp 1644511149
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_317
timestamp 1644511149
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1644511149
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1644511149
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_337
timestamp 1644511149
transform 1 0 32108 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_345
timestamp 1644511149
transform 1 0 32844 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_367
timestamp 1644511149
transform 1 0 34868 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_379
timestamp 1644511149
transform 1 0 35972 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1644511149
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_393
timestamp 1644511149
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_405
timestamp 1644511149
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_417
timestamp 1644511149
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_429
timestamp 1644511149
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1644511149
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1644511149
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_449
timestamp 1644511149
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_461
timestamp 1644511149
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_473
timestamp 1644511149
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_485
timestamp 1644511149
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1644511149
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1644511149
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_505
timestamp 1644511149
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_517
timestamp 1644511149
transform 1 0 48668 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_544
timestamp 1644511149
transform 1 0 51152 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_556
timestamp 1644511149
transform 1 0 52256 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_561
timestamp 1644511149
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_573
timestamp 1644511149
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_585
timestamp 1644511149
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_597
timestamp 1644511149
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1644511149
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1644511149
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_617
timestamp 1644511149
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_629
timestamp 1644511149
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_641
timestamp 1644511149
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_653
timestamp 1644511149
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_665
timestamp 1644511149
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1644511149
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_673
timestamp 1644511149
transform 1 0 63020 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_681
timestamp 1644511149
transform 1 0 63756 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_704
timestamp 1644511149
transform 1 0 65872 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_716
timestamp 1644511149
transform 1 0 66976 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_729
timestamp 1644511149
transform 1 0 68172 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_3
timestamp 1644511149
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_15
timestamp 1644511149
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1644511149
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_29
timestamp 1644511149
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_41
timestamp 1644511149
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_53
timestamp 1644511149
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_65
timestamp 1644511149
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1644511149
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1644511149
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_85
timestamp 1644511149
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_97
timestamp 1644511149
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_109
timestamp 1644511149
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_121
timestamp 1644511149
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1644511149
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1644511149
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_141
timestamp 1644511149
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_153
timestamp 1644511149
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_165
timestamp 1644511149
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_177
timestamp 1644511149
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1644511149
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1644511149
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_197
timestamp 1644511149
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_209
timestamp 1644511149
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_221
timestamp 1644511149
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_233
timestamp 1644511149
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1644511149
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1644511149
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_253
timestamp 1644511149
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_265
timestamp 1644511149
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_277
timestamp 1644511149
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_289
timestamp 1644511149
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1644511149
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1644511149
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_309
timestamp 1644511149
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_321
timestamp 1644511149
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_333
timestamp 1644511149
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_345
timestamp 1644511149
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1644511149
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1644511149
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_368
timestamp 1644511149
transform 1 0 34960 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_380
timestamp 1644511149
transform 1 0 36064 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_392
timestamp 1644511149
transform 1 0 37168 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_404
timestamp 1644511149
transform 1 0 38272 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_416
timestamp 1644511149
transform 1 0 39376 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_421
timestamp 1644511149
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_433
timestamp 1644511149
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_445
timestamp 1644511149
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_457
timestamp 1644511149
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1644511149
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1644511149
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_477
timestamp 1644511149
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_489
timestamp 1644511149
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_501
timestamp 1644511149
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_513
timestamp 1644511149
transform 1 0 48300 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_521
timestamp 1644511149
transform 1 0 49036 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_100_526
timestamp 1644511149
transform 1 0 49496 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_100_533
timestamp 1644511149
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_545
timestamp 1644511149
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_557
timestamp 1644511149
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_569
timestamp 1644511149
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1644511149
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1644511149
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_589
timestamp 1644511149
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_601
timestamp 1644511149
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_613
timestamp 1644511149
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_625
timestamp 1644511149
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_637
timestamp 1644511149
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_643
timestamp 1644511149
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_645
timestamp 1644511149
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_657
timestamp 1644511149
transform 1 0 61548 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_669
timestamp 1644511149
transform 1 0 62652 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_681
timestamp 1644511149
transform 1 0 63756 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_687
timestamp 1644511149
transform 1 0 64308 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_699
timestamp 1644511149
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_701
timestamp 1644511149
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_713
timestamp 1644511149
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_725
timestamp 1644511149
transform 1 0 67804 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1644511149
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1644511149
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_27
timestamp 1644511149
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_39
timestamp 1644511149
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1644511149
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1644511149
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1644511149
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1644511149
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_81
timestamp 1644511149
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_93
timestamp 1644511149
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1644511149
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1644511149
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_113
timestamp 1644511149
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_125
timestamp 1644511149
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_137
timestamp 1644511149
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_149
timestamp 1644511149
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_161
timestamp 1644511149
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1644511149
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_169
timestamp 1644511149
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_181
timestamp 1644511149
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_193
timestamp 1644511149
transform 1 0 18860 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_205
timestamp 1644511149
transform 1 0 19964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_217
timestamp 1644511149
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1644511149
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_225
timestamp 1644511149
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_237
timestamp 1644511149
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_249
timestamp 1644511149
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_261
timestamp 1644511149
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1644511149
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1644511149
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_281
timestamp 1644511149
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_293
timestamp 1644511149
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_305
timestamp 1644511149
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_317
timestamp 1644511149
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_329
timestamp 1644511149
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_335
timestamp 1644511149
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_337
timestamp 1644511149
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_349
timestamp 1644511149
transform 1 0 33212 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_357
timestamp 1644511149
transform 1 0 33948 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_381
timestamp 1644511149
transform 1 0 36156 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 1644511149
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_393
timestamp 1644511149
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_405
timestamp 1644511149
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_417
timestamp 1644511149
transform 1 0 39468 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_429
timestamp 1644511149
transform 1 0 40572 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1644511149
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1644511149
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_449
timestamp 1644511149
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_461
timestamp 1644511149
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_473
timestamp 1644511149
transform 1 0 44620 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_485
timestamp 1644511149
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1644511149
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1644511149
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_505
timestamp 1644511149
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_517
timestamp 1644511149
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_529
timestamp 1644511149
transform 1 0 49772 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_541
timestamp 1644511149
transform 1 0 50876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_553
timestamp 1644511149
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1644511149
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_561
timestamp 1644511149
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_573
timestamp 1644511149
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_585
timestamp 1644511149
transform 1 0 54924 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_597
timestamp 1644511149
transform 1 0 56028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_609
timestamp 1644511149
transform 1 0 57132 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1644511149
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_617
timestamp 1644511149
transform 1 0 57868 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_629
timestamp 1644511149
transform 1 0 58972 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_641
timestamp 1644511149
transform 1 0 60076 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_653
timestamp 1644511149
transform 1 0 61180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_665
timestamp 1644511149
transform 1 0 62284 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_671
timestamp 1644511149
transform 1 0 62836 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_673
timestamp 1644511149
transform 1 0 63020 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_681
timestamp 1644511149
transform 1 0 63756 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_705
timestamp 1644511149
transform 1 0 65964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_717
timestamp 1644511149
transform 1 0 67068 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_725
timestamp 1644511149
transform 1 0 67804 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_729
timestamp 1644511149
transform 1 0 68172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_3
timestamp 1644511149
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_15
timestamp 1644511149
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1644511149
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_29
timestamp 1644511149
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_41
timestamp 1644511149
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_53
timestamp 1644511149
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1644511149
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1644511149
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1644511149
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_85
timestamp 1644511149
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_97
timestamp 1644511149
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_109
timestamp 1644511149
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_121
timestamp 1644511149
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1644511149
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1644511149
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_141
timestamp 1644511149
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_153
timestamp 1644511149
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_165
timestamp 1644511149
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_177
timestamp 1644511149
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_189
timestamp 1644511149
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1644511149
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_197
timestamp 1644511149
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_209
timestamp 1644511149
transform 1 0 20332 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_221
timestamp 1644511149
transform 1 0 21436 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_233
timestamp 1644511149
transform 1 0 22540 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_245
timestamp 1644511149
transform 1 0 23644 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_251
timestamp 1644511149
transform 1 0 24196 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_253
timestamp 1644511149
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_265
timestamp 1644511149
transform 1 0 25484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_277
timestamp 1644511149
transform 1 0 26588 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_289
timestamp 1644511149
transform 1 0 27692 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_301
timestamp 1644511149
transform 1 0 28796 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_307
timestamp 1644511149
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_309
timestamp 1644511149
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_321
timestamp 1644511149
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_333
timestamp 1644511149
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_345
timestamp 1644511149
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_357
timestamp 1644511149
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_363
timestamp 1644511149
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_368
timestamp 1644511149
transform 1 0 34960 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_380
timestamp 1644511149
transform 1 0 36064 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_102_403
timestamp 1644511149
transform 1 0 38180 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_415
timestamp 1644511149
transform 1 0 39284 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_419
timestamp 1644511149
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_421
timestamp 1644511149
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_433
timestamp 1644511149
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_445
timestamp 1644511149
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_457
timestamp 1644511149
transform 1 0 43148 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_469
timestamp 1644511149
transform 1 0 44252 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_475
timestamp 1644511149
transform 1 0 44804 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_477
timestamp 1644511149
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_489
timestamp 1644511149
transform 1 0 46092 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_501
timestamp 1644511149
transform 1 0 47196 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_513
timestamp 1644511149
transform 1 0 48300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_525
timestamp 1644511149
transform 1 0 49404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_531
timestamp 1644511149
transform 1 0 49956 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_533
timestamp 1644511149
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_545
timestamp 1644511149
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_557
timestamp 1644511149
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_569
timestamp 1644511149
transform 1 0 53452 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_581
timestamp 1644511149
transform 1 0 54556 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_587
timestamp 1644511149
transform 1 0 55108 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_589
timestamp 1644511149
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_601
timestamp 1644511149
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_613
timestamp 1644511149
transform 1 0 57500 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_625
timestamp 1644511149
transform 1 0 58604 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_637
timestamp 1644511149
transform 1 0 59708 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_643
timestamp 1644511149
transform 1 0 60260 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_645
timestamp 1644511149
transform 1 0 60444 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_657
timestamp 1644511149
transform 1 0 61548 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_669
timestamp 1644511149
transform 1 0 62652 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_675
timestamp 1644511149
transform 1 0 63204 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_679
timestamp 1644511149
transform 1 0 63572 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_686
timestamp 1644511149
transform 1 0 64216 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_102_693
timestamp 1644511149
transform 1 0 64860 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_699
timestamp 1644511149
transform 1 0 65412 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_704
timestamp 1644511149
transform 1 0 65872 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_716
timestamp 1644511149
transform 1 0 66976 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_728
timestamp 1644511149
transform 1 0 68080 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_732
timestamp 1644511149
transform 1 0 68448 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_3
timestamp 1644511149
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_15
timestamp 1644511149
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_27
timestamp 1644511149
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_39
timestamp 1644511149
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_51
timestamp 1644511149
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1644511149
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1644511149
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1644511149
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_81
timestamp 1644511149
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_93
timestamp 1644511149
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1644511149
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1644511149
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_113
timestamp 1644511149
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_125
timestamp 1644511149
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_137
timestamp 1644511149
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_149
timestamp 1644511149
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_161
timestamp 1644511149
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_167
timestamp 1644511149
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_169
timestamp 1644511149
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_181
timestamp 1644511149
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_193
timestamp 1644511149
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_205
timestamp 1644511149
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_217
timestamp 1644511149
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_223
timestamp 1644511149
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_225
timestamp 1644511149
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_237
timestamp 1644511149
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_249
timestamp 1644511149
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_261
timestamp 1644511149
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_273
timestamp 1644511149
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_279
timestamp 1644511149
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_281
timestamp 1644511149
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_293
timestamp 1644511149
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_305
timestamp 1644511149
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_317
timestamp 1644511149
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_329
timestamp 1644511149
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_335
timestamp 1644511149
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_337
timestamp 1644511149
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_349
timestamp 1644511149
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_361
timestamp 1644511149
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_373
timestamp 1644511149
transform 1 0 35420 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_378
timestamp 1644511149
transform 1 0 35880 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_382
timestamp 1644511149
transform 1 0 36248 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_103_386
timestamp 1644511149
transform 1 0 36616 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_103_396
timestamp 1644511149
transform 1 0 37536 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_408
timestamp 1644511149
transform 1 0 38640 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_420
timestamp 1644511149
transform 1 0 39744 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_432
timestamp 1644511149
transform 1 0 40848 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_444
timestamp 1644511149
transform 1 0 41952 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_449
timestamp 1644511149
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_461
timestamp 1644511149
transform 1 0 43516 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_473
timestamp 1644511149
transform 1 0 44620 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_485
timestamp 1644511149
transform 1 0 45724 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_497
timestamp 1644511149
transform 1 0 46828 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_503
timestamp 1644511149
transform 1 0 47380 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_505
timestamp 1644511149
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_517
timestamp 1644511149
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_529
timestamp 1644511149
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_541
timestamp 1644511149
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_553
timestamp 1644511149
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_559
timestamp 1644511149
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_561
timestamp 1644511149
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_573
timestamp 1644511149
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_585
timestamp 1644511149
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_597
timestamp 1644511149
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_609
timestamp 1644511149
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_615
timestamp 1644511149
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_617
timestamp 1644511149
transform 1 0 57868 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_629
timestamp 1644511149
transform 1 0 58972 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_641
timestamp 1644511149
transform 1 0 60076 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_653
timestamp 1644511149
transform 1 0 61180 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_665
timestamp 1644511149
transform 1 0 62284 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_671
timestamp 1644511149
transform 1 0 62836 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_673
timestamp 1644511149
transform 1 0 63020 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_685
timestamp 1644511149
transform 1 0 64124 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_103_708
timestamp 1644511149
transform 1 0 66240 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_720
timestamp 1644511149
transform 1 0 67344 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_103_729
timestamp 1644511149
transform 1 0 68172 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_3
timestamp 1644511149
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_15
timestamp 1644511149
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1644511149
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1644511149
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_41
timestamp 1644511149
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_53
timestamp 1644511149
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_65
timestamp 1644511149
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1644511149
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1644511149
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_85
timestamp 1644511149
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_97
timestamp 1644511149
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_109
timestamp 1644511149
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_121
timestamp 1644511149
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1644511149
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1644511149
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_141
timestamp 1644511149
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_153
timestamp 1644511149
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_165
timestamp 1644511149
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_177
timestamp 1644511149
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_189
timestamp 1644511149
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_195
timestamp 1644511149
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_197
timestamp 1644511149
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_209
timestamp 1644511149
transform 1 0 20332 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_221
timestamp 1644511149
transform 1 0 21436 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_233
timestamp 1644511149
transform 1 0 22540 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_245
timestamp 1644511149
transform 1 0 23644 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_251
timestamp 1644511149
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_253
timestamp 1644511149
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_265
timestamp 1644511149
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_277
timestamp 1644511149
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_289
timestamp 1644511149
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_301
timestamp 1644511149
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_307
timestamp 1644511149
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_309
timestamp 1644511149
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_321
timestamp 1644511149
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_333
timestamp 1644511149
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_345
timestamp 1644511149
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_357
timestamp 1644511149
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_363
timestamp 1644511149
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_365
timestamp 1644511149
transform 1 0 34684 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_373
timestamp 1644511149
transform 1 0 35420 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_395
timestamp 1644511149
transform 1 0 37444 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_407
timestamp 1644511149
transform 1 0 38548 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_419
timestamp 1644511149
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_421
timestamp 1644511149
transform 1 0 39836 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_433
timestamp 1644511149
transform 1 0 40940 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_445
timestamp 1644511149
transform 1 0 42044 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_457
timestamp 1644511149
transform 1 0 43148 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_469
timestamp 1644511149
transform 1 0 44252 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_475
timestamp 1644511149
transform 1 0 44804 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_477
timestamp 1644511149
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_489
timestamp 1644511149
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_501
timestamp 1644511149
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_513
timestamp 1644511149
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_525
timestamp 1644511149
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_531
timestamp 1644511149
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_533
timestamp 1644511149
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_545
timestamp 1644511149
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_557
timestamp 1644511149
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_569
timestamp 1644511149
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_581
timestamp 1644511149
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_587
timestamp 1644511149
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_589
timestamp 1644511149
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_601
timestamp 1644511149
transform 1 0 56396 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_613
timestamp 1644511149
transform 1 0 57500 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_625
timestamp 1644511149
transform 1 0 58604 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_637
timestamp 1644511149
transform 1 0 59708 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_643
timestamp 1644511149
transform 1 0 60260 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_645
timestamp 1644511149
transform 1 0 60444 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_657
timestamp 1644511149
transform 1 0 61548 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_669
timestamp 1644511149
transform 1 0 62652 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_681
timestamp 1644511149
transform 1 0 63756 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_693
timestamp 1644511149
transform 1 0 64860 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_699
timestamp 1644511149
transform 1 0 65412 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_701
timestamp 1644511149
transform 1 0 65596 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_713
timestamp 1644511149
transform 1 0 66700 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_725
timestamp 1644511149
transform 1 0 67804 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_3
timestamp 1644511149
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1644511149
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1644511149
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_39
timestamp 1644511149
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1644511149
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1644511149
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1644511149
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1644511149
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_81
timestamp 1644511149
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_93
timestamp 1644511149
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1644511149
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1644511149
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_113
timestamp 1644511149
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_125
timestamp 1644511149
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_137
timestamp 1644511149
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_149
timestamp 1644511149
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1644511149
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1644511149
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_169
timestamp 1644511149
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_181
timestamp 1644511149
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_193
timestamp 1644511149
transform 1 0 18860 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_205
timestamp 1644511149
transform 1 0 19964 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_217
timestamp 1644511149
transform 1 0 21068 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_223
timestamp 1644511149
transform 1 0 21620 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_225
timestamp 1644511149
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_237
timestamp 1644511149
transform 1 0 22908 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_249
timestamp 1644511149
transform 1 0 24012 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_261
timestamp 1644511149
transform 1 0 25116 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_276
timestamp 1644511149
transform 1 0 26496 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_302
timestamp 1644511149
transform 1 0 28888 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_314
timestamp 1644511149
transform 1 0 29992 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_326
timestamp 1644511149
transform 1 0 31096 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_334
timestamp 1644511149
transform 1 0 31832 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_337
timestamp 1644511149
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_349
timestamp 1644511149
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_361
timestamp 1644511149
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_373
timestamp 1644511149
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_385
timestamp 1644511149
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_391
timestamp 1644511149
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_393
timestamp 1644511149
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_405
timestamp 1644511149
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_417
timestamp 1644511149
transform 1 0 39468 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_429
timestamp 1644511149
transform 1 0 40572 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_441
timestamp 1644511149
transform 1 0 41676 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_447
timestamp 1644511149
transform 1 0 42228 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_449
timestamp 1644511149
transform 1 0 42412 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_461
timestamp 1644511149
transform 1 0 43516 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_473
timestamp 1644511149
transform 1 0 44620 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_485
timestamp 1644511149
transform 1 0 45724 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_497
timestamp 1644511149
transform 1 0 46828 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_503
timestamp 1644511149
transform 1 0 47380 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_505
timestamp 1644511149
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_517
timestamp 1644511149
transform 1 0 48668 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_529
timestamp 1644511149
transform 1 0 49772 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_541
timestamp 1644511149
transform 1 0 50876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_553
timestamp 1644511149
transform 1 0 51980 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_559
timestamp 1644511149
transform 1 0 52532 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_561
timestamp 1644511149
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_573
timestamp 1644511149
transform 1 0 53820 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_580
timestamp 1644511149
transform 1 0 54464 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_105_605
timestamp 1644511149
transform 1 0 56764 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_105_613
timestamp 1644511149
transform 1 0 57500 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_617
timestamp 1644511149
transform 1 0 57868 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_629
timestamp 1644511149
transform 1 0 58972 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_641
timestamp 1644511149
transform 1 0 60076 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_653
timestamp 1644511149
transform 1 0 61180 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_665
timestamp 1644511149
transform 1 0 62284 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_671
timestamp 1644511149
transform 1 0 62836 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_673
timestamp 1644511149
transform 1 0 63020 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_685
timestamp 1644511149
transform 1 0 64124 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_697
timestamp 1644511149
transform 1 0 65228 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_709
timestamp 1644511149
transform 1 0 66332 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_721
timestamp 1644511149
transform 1 0 67436 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_727
timestamp 1644511149
transform 1 0 67988 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_729
timestamp 1644511149
transform 1 0 68172 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_3
timestamp 1644511149
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_15
timestamp 1644511149
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1644511149
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1644511149
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1644511149
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1644511149
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_65
timestamp 1644511149
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1644511149
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1644511149
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_85
timestamp 1644511149
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_97
timestamp 1644511149
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_109
timestamp 1644511149
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_121
timestamp 1644511149
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_133
timestamp 1644511149
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1644511149
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_141
timestamp 1644511149
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_153
timestamp 1644511149
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_165
timestamp 1644511149
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_177
timestamp 1644511149
transform 1 0 17388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_189
timestamp 1644511149
transform 1 0 18492 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_195
timestamp 1644511149
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_197
timestamp 1644511149
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_209
timestamp 1644511149
transform 1 0 20332 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_221
timestamp 1644511149
transform 1 0 21436 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_233
timestamp 1644511149
transform 1 0 22540 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_245
timestamp 1644511149
transform 1 0 23644 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_251
timestamp 1644511149
transform 1 0 24196 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_253
timestamp 1644511149
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_265
timestamp 1644511149
transform 1 0 25484 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_273
timestamp 1644511149
transform 1 0 26220 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_277
timestamp 1644511149
transform 1 0 26588 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_289
timestamp 1644511149
transform 1 0 27692 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_301
timestamp 1644511149
transform 1 0 28796 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_307
timestamp 1644511149
transform 1 0 29348 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_309
timestamp 1644511149
transform 1 0 29532 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_321
timestamp 1644511149
transform 1 0 30636 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_333
timestamp 1644511149
transform 1 0 31740 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_345
timestamp 1644511149
transform 1 0 32844 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_357
timestamp 1644511149
transform 1 0 33948 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_363
timestamp 1644511149
transform 1 0 34500 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_365
timestamp 1644511149
transform 1 0 34684 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_373
timestamp 1644511149
transform 1 0 35420 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_106_378
timestamp 1644511149
transform 1 0 35880 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_390
timestamp 1644511149
transform 1 0 36984 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_402
timestamp 1644511149
transform 1 0 38088 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_414
timestamp 1644511149
transform 1 0 39192 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_106_421
timestamp 1644511149
transform 1 0 39836 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_433
timestamp 1644511149
transform 1 0 40940 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_445
timestamp 1644511149
transform 1 0 42044 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_457
timestamp 1644511149
transform 1 0 43148 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_469
timestamp 1644511149
transform 1 0 44252 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_475
timestamp 1644511149
transform 1 0 44804 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_477
timestamp 1644511149
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_489
timestamp 1644511149
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_501
timestamp 1644511149
transform 1 0 47196 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_513
timestamp 1644511149
transform 1 0 48300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_525
timestamp 1644511149
transform 1 0 49404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1644511149
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_533
timestamp 1644511149
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_545
timestamp 1644511149
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_557
timestamp 1644511149
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_569
timestamp 1644511149
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_581
timestamp 1644511149
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_587
timestamp 1644511149
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_592
timestamp 1644511149
transform 1 0 55568 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_604
timestamp 1644511149
transform 1 0 56672 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_616
timestamp 1644511149
transform 1 0 57776 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_628
timestamp 1644511149
transform 1 0 58880 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_640
timestamp 1644511149
transform 1 0 59984 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_645
timestamp 1644511149
transform 1 0 60444 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_657
timestamp 1644511149
transform 1 0 61548 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_669
timestamp 1644511149
transform 1 0 62652 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_681
timestamp 1644511149
transform 1 0 63756 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_693
timestamp 1644511149
transform 1 0 64860 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_699
timestamp 1644511149
transform 1 0 65412 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_701
timestamp 1644511149
transform 1 0 65596 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_713
timestamp 1644511149
transform 1 0 66700 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_725
timestamp 1644511149
transform 1 0 67804 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_3
timestamp 1644511149
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_15
timestamp 1644511149
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_27
timestamp 1644511149
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_39
timestamp 1644511149
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_51
timestamp 1644511149
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1644511149
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1644511149
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1644511149
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_81
timestamp 1644511149
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_93
timestamp 1644511149
transform 1 0 9660 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_105
timestamp 1644511149
transform 1 0 10764 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_111
timestamp 1644511149
transform 1 0 11316 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_113
timestamp 1644511149
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_125
timestamp 1644511149
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_137
timestamp 1644511149
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_149
timestamp 1644511149
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_161
timestamp 1644511149
transform 1 0 15916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_167
timestamp 1644511149
transform 1 0 16468 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_169
timestamp 1644511149
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_181
timestamp 1644511149
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_193
timestamp 1644511149
transform 1 0 18860 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_205
timestamp 1644511149
transform 1 0 19964 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_217
timestamp 1644511149
transform 1 0 21068 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_223
timestamp 1644511149
transform 1 0 21620 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_225
timestamp 1644511149
transform 1 0 21804 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_237
timestamp 1644511149
transform 1 0 22908 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_249
timestamp 1644511149
transform 1 0 24012 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_261
timestamp 1644511149
transform 1 0 25116 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_273
timestamp 1644511149
transform 1 0 26220 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_279
timestamp 1644511149
transform 1 0 26772 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_281
timestamp 1644511149
transform 1 0 26956 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_293
timestamp 1644511149
transform 1 0 28060 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_305
timestamp 1644511149
transform 1 0 29164 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_317
timestamp 1644511149
transform 1 0 30268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_329
timestamp 1644511149
transform 1 0 31372 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_335
timestamp 1644511149
transform 1 0 31924 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_337
timestamp 1644511149
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_349
timestamp 1644511149
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_361
timestamp 1644511149
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_373
timestamp 1644511149
transform 1 0 35420 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_385
timestamp 1644511149
transform 1 0 36524 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_391
timestamp 1644511149
transform 1 0 37076 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_393
timestamp 1644511149
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_405
timestamp 1644511149
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_417
timestamp 1644511149
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_429
timestamp 1644511149
transform 1 0 40572 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_441
timestamp 1644511149
transform 1 0 41676 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_447
timestamp 1644511149
transform 1 0 42228 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_449
timestamp 1644511149
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_461
timestamp 1644511149
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_473
timestamp 1644511149
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_485
timestamp 1644511149
transform 1 0 45724 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_107_490
timestamp 1644511149
transform 1 0 46184 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_502
timestamp 1644511149
transform 1 0 47288 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_107_505
timestamp 1644511149
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_517
timestamp 1644511149
transform 1 0 48668 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_529
timestamp 1644511149
transform 1 0 49772 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_541
timestamp 1644511149
transform 1 0 50876 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_553
timestamp 1644511149
transform 1 0 51980 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_559
timestamp 1644511149
transform 1 0 52532 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_561
timestamp 1644511149
transform 1 0 52716 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_573
timestamp 1644511149
transform 1 0 53820 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_585
timestamp 1644511149
transform 1 0 54924 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_597
timestamp 1644511149
transform 1 0 56028 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_609
timestamp 1644511149
transform 1 0 57132 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_615
timestamp 1644511149
transform 1 0 57684 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_617
timestamp 1644511149
transform 1 0 57868 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_629
timestamp 1644511149
transform 1 0 58972 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_641
timestamp 1644511149
transform 1 0 60076 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_653
timestamp 1644511149
transform 1 0 61180 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_665
timestamp 1644511149
transform 1 0 62284 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_671
timestamp 1644511149
transform 1 0 62836 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_673
timestamp 1644511149
transform 1 0 63020 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_685
timestamp 1644511149
transform 1 0 64124 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_697
timestamp 1644511149
transform 1 0 65228 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_709
timestamp 1644511149
transform 1 0 66332 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_721
timestamp 1644511149
transform 1 0 67436 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_727
timestamp 1644511149
transform 1 0 67988 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_729
timestamp 1644511149
transform 1 0 68172 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_108_3
timestamp 1644511149
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_15
timestamp 1644511149
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1644511149
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_29
timestamp 1644511149
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_41
timestamp 1644511149
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_53
timestamp 1644511149
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_65
timestamp 1644511149
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1644511149
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1644511149
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_85
timestamp 1644511149
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_97
timestamp 1644511149
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_109
timestamp 1644511149
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_121
timestamp 1644511149
transform 1 0 12236 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_133
timestamp 1644511149
transform 1 0 13340 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_139
timestamp 1644511149
transform 1 0 13892 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_141
timestamp 1644511149
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_153
timestamp 1644511149
transform 1 0 15180 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_165
timestamp 1644511149
transform 1 0 16284 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_177
timestamp 1644511149
transform 1 0 17388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_189
timestamp 1644511149
transform 1 0 18492 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_195
timestamp 1644511149
transform 1 0 19044 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_197
timestamp 1644511149
transform 1 0 19228 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_209
timestamp 1644511149
transform 1 0 20332 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_221
timestamp 1644511149
transform 1 0 21436 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_233
timestamp 1644511149
transform 1 0 22540 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_245
timestamp 1644511149
transform 1 0 23644 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_251
timestamp 1644511149
transform 1 0 24196 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_253
timestamp 1644511149
transform 1 0 24380 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_265
timestamp 1644511149
transform 1 0 25484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_277
timestamp 1644511149
transform 1 0 26588 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_289
timestamp 1644511149
transform 1 0 27692 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_301
timestamp 1644511149
transform 1 0 28796 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_307
timestamp 1644511149
transform 1 0 29348 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_309
timestamp 1644511149
transform 1 0 29532 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_321
timestamp 1644511149
transform 1 0 30636 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_333
timestamp 1644511149
transform 1 0 31740 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_345
timestamp 1644511149
transform 1 0 32844 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_357
timestamp 1644511149
transform 1 0 33948 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_363
timestamp 1644511149
transform 1 0 34500 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_365
timestamp 1644511149
transform 1 0 34684 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_377
timestamp 1644511149
transform 1 0 35788 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_389
timestamp 1644511149
transform 1 0 36892 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_401
timestamp 1644511149
transform 1 0 37996 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_413
timestamp 1644511149
transform 1 0 39100 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_419
timestamp 1644511149
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_421
timestamp 1644511149
transform 1 0 39836 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_433
timestamp 1644511149
transform 1 0 40940 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_445
timestamp 1644511149
transform 1 0 42044 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_457
timestamp 1644511149
transform 1 0 43148 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_469
timestamp 1644511149
transform 1 0 44252 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_475
timestamp 1644511149
transform 1 0 44804 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_477
timestamp 1644511149
transform 1 0 44988 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_485
timestamp 1644511149
transform 1 0 45724 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_507
timestamp 1644511149
transform 1 0 47748 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_519
timestamp 1644511149
transform 1 0 48852 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1644511149
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_533
timestamp 1644511149
transform 1 0 50140 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_545
timestamp 1644511149
transform 1 0 51244 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_557
timestamp 1644511149
transform 1 0 52348 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_569
timestamp 1644511149
transform 1 0 53452 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_575
timestamp 1644511149
transform 1 0 54004 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_579
timestamp 1644511149
transform 1 0 54372 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_587
timestamp 1644511149
transform 1 0 55108 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_610
timestamp 1644511149
transform 1 0 57224 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_622
timestamp 1644511149
transform 1 0 58328 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_634
timestamp 1644511149
transform 1 0 59432 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_642
timestamp 1644511149
transform 1 0 60168 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_108_645
timestamp 1644511149
transform 1 0 60444 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_657
timestamp 1644511149
transform 1 0 61548 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_669
timestamp 1644511149
transform 1 0 62652 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_681
timestamp 1644511149
transform 1 0 63756 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_693
timestamp 1644511149
transform 1 0 64860 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_699
timestamp 1644511149
transform 1 0 65412 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_701
timestamp 1644511149
transform 1 0 65596 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_713
timestamp 1644511149
transform 1 0 66700 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_725
timestamp 1644511149
transform 1 0 67804 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_3
timestamp 1644511149
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_15
timestamp 1644511149
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_27
timestamp 1644511149
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_39
timestamp 1644511149
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1644511149
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1644511149
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1644511149
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1644511149
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_81
timestamp 1644511149
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_93
timestamp 1644511149
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_105
timestamp 1644511149
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_111
timestamp 1644511149
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_113
timestamp 1644511149
transform 1 0 11500 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_125
timestamp 1644511149
transform 1 0 12604 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_137
timestamp 1644511149
transform 1 0 13708 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_149
timestamp 1644511149
transform 1 0 14812 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_161
timestamp 1644511149
transform 1 0 15916 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_167
timestamp 1644511149
transform 1 0 16468 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_169
timestamp 1644511149
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_181
timestamp 1644511149
transform 1 0 17756 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_193
timestamp 1644511149
transform 1 0 18860 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_205
timestamp 1644511149
transform 1 0 19964 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_217
timestamp 1644511149
transform 1 0 21068 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_223
timestamp 1644511149
transform 1 0 21620 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_225
timestamp 1644511149
transform 1 0 21804 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_237
timestamp 1644511149
transform 1 0 22908 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_249
timestamp 1644511149
transform 1 0 24012 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_261
timestamp 1644511149
transform 1 0 25116 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_273
timestamp 1644511149
transform 1 0 26220 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_279
timestamp 1644511149
transform 1 0 26772 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_281
timestamp 1644511149
transform 1 0 26956 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_293
timestamp 1644511149
transform 1 0 28060 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_305
timestamp 1644511149
transform 1 0 29164 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_317
timestamp 1644511149
transform 1 0 30268 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_109_328
timestamp 1644511149
transform 1 0 31280 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_340
timestamp 1644511149
transform 1 0 32384 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_352
timestamp 1644511149
transform 1 0 33488 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_364
timestamp 1644511149
transform 1 0 34592 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_376
timestamp 1644511149
transform 1 0 35696 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_109_384
timestamp 1644511149
transform 1 0 36432 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_109_388
timestamp 1644511149
transform 1 0 36800 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_109_414
timestamp 1644511149
transform 1 0 39192 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_426
timestamp 1644511149
transform 1 0 40296 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_438
timestamp 1644511149
transform 1 0 41400 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_446
timestamp 1644511149
transform 1 0 42136 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_449
timestamp 1644511149
transform 1 0 42412 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_461
timestamp 1644511149
transform 1 0 43516 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_473
timestamp 1644511149
transform 1 0 44620 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_485
timestamp 1644511149
transform 1 0 45724 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_490
timestamp 1644511149
transform 1 0 46184 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_502
timestamp 1644511149
transform 1 0 47288 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_505
timestamp 1644511149
transform 1 0 47564 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_517
timestamp 1644511149
transform 1 0 48668 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_529
timestamp 1644511149
transform 1 0 49772 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_541
timestamp 1644511149
transform 1 0 50876 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_553
timestamp 1644511149
transform 1 0 51980 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_559
timestamp 1644511149
transform 1 0 52532 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_561
timestamp 1644511149
transform 1 0 52716 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_573
timestamp 1644511149
transform 1 0 53820 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_584
timestamp 1644511149
transform 1 0 54832 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_596
timestamp 1644511149
transform 1 0 55936 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_608
timestamp 1644511149
transform 1 0 57040 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_617
timestamp 1644511149
transform 1 0 57868 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_629
timestamp 1644511149
transform 1 0 58972 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_641
timestamp 1644511149
transform 1 0 60076 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_653
timestamp 1644511149
transform 1 0 61180 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_665
timestamp 1644511149
transform 1 0 62284 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_671
timestamp 1644511149
transform 1 0 62836 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_673
timestamp 1644511149
transform 1 0 63020 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_685
timestamp 1644511149
transform 1 0 64124 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_697
timestamp 1644511149
transform 1 0 65228 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_709
timestamp 1644511149
transform 1 0 66332 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_721
timestamp 1644511149
transform 1 0 67436 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_727
timestamp 1644511149
transform 1 0 67988 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_109_729
timestamp 1644511149
transform 1 0 68172 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_110_3
timestamp 1644511149
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_15
timestamp 1644511149
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1644511149
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1644511149
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1644511149
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1644511149
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_65
timestamp 1644511149
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1644511149
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1644511149
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_85
timestamp 1644511149
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_97
timestamp 1644511149
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_109
timestamp 1644511149
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_121
timestamp 1644511149
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_133
timestamp 1644511149
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_139
timestamp 1644511149
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_141
timestamp 1644511149
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_153
timestamp 1644511149
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_165
timestamp 1644511149
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_177
timestamp 1644511149
transform 1 0 17388 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_189
timestamp 1644511149
transform 1 0 18492 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_195
timestamp 1644511149
transform 1 0 19044 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_197
timestamp 1644511149
transform 1 0 19228 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_209
timestamp 1644511149
transform 1 0 20332 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_221
timestamp 1644511149
transform 1 0 21436 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_233
timestamp 1644511149
transform 1 0 22540 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_245
timestamp 1644511149
transform 1 0 23644 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_251
timestamp 1644511149
transform 1 0 24196 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_253
timestamp 1644511149
transform 1 0 24380 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_265
timestamp 1644511149
transform 1 0 25484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_277
timestamp 1644511149
transform 1 0 26588 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_289
timestamp 1644511149
transform 1 0 27692 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_301
timestamp 1644511149
transform 1 0 28796 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_307
timestamp 1644511149
transform 1 0 29348 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_309
timestamp 1644511149
transform 1 0 29532 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_110_321
timestamp 1644511149
transform 1 0 30636 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_345
timestamp 1644511149
transform 1 0 32844 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_357
timestamp 1644511149
transform 1 0 33948 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_363
timestamp 1644511149
transform 1 0 34500 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_365
timestamp 1644511149
transform 1 0 34684 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_377
timestamp 1644511149
transform 1 0 35788 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_392
timestamp 1644511149
transform 1 0 37168 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_404
timestamp 1644511149
transform 1 0 38272 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_416
timestamp 1644511149
transform 1 0 39376 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_110_421
timestamp 1644511149
transform 1 0 39836 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_433
timestamp 1644511149
transform 1 0 40940 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_445
timestamp 1644511149
transform 1 0 42044 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_457
timestamp 1644511149
transform 1 0 43148 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_469
timestamp 1644511149
transform 1 0 44252 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_475
timestamp 1644511149
transform 1 0 44804 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_477
timestamp 1644511149
transform 1 0 44988 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_489
timestamp 1644511149
transform 1 0 46092 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_501
timestamp 1644511149
transform 1 0 47196 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_513
timestamp 1644511149
transform 1 0 48300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_525
timestamp 1644511149
transform 1 0 49404 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_531
timestamp 1644511149
transform 1 0 49956 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_533
timestamp 1644511149
transform 1 0 50140 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_545
timestamp 1644511149
transform 1 0 51244 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_557
timestamp 1644511149
transform 1 0 52348 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_569
timestamp 1644511149
transform 1 0 53452 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_581
timestamp 1644511149
transform 1 0 54556 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_587
timestamp 1644511149
transform 1 0 55108 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_589
timestamp 1644511149
transform 1 0 55292 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_601
timestamp 1644511149
transform 1 0 56396 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_613
timestamp 1644511149
transform 1 0 57500 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_625
timestamp 1644511149
transform 1 0 58604 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_637
timestamp 1644511149
transform 1 0 59708 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_643
timestamp 1644511149
transform 1 0 60260 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_645
timestamp 1644511149
transform 1 0 60444 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_657
timestamp 1644511149
transform 1 0 61548 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_669
timestamp 1644511149
transform 1 0 62652 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_681
timestamp 1644511149
transform 1 0 63756 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_693
timestamp 1644511149
transform 1 0 64860 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_699
timestamp 1644511149
transform 1 0 65412 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_701
timestamp 1644511149
transform 1 0 65596 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_713
timestamp 1644511149
transform 1 0 66700 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_725
timestamp 1644511149
transform 1 0 67804 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_3
timestamp 1644511149
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_15
timestamp 1644511149
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_27
timestamp 1644511149
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_39
timestamp 1644511149
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1644511149
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1644511149
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_57
timestamp 1644511149
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_69
timestamp 1644511149
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_81
timestamp 1644511149
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_93
timestamp 1644511149
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_105
timestamp 1644511149
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_111
timestamp 1644511149
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_113
timestamp 1644511149
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_125
timestamp 1644511149
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_137
timestamp 1644511149
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_149
timestamp 1644511149
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_161
timestamp 1644511149
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_167
timestamp 1644511149
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_169
timestamp 1644511149
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_181
timestamp 1644511149
transform 1 0 17756 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_193
timestamp 1644511149
transform 1 0 18860 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_111_202
timestamp 1644511149
transform 1 0 19688 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_209
timestamp 1644511149
transform 1 0 20332 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_221
timestamp 1644511149
transform 1 0 21436 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_111_225
timestamp 1644511149
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_237
timestamp 1644511149
transform 1 0 22908 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_249
timestamp 1644511149
transform 1 0 24012 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_261
timestamp 1644511149
transform 1 0 25116 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_273
timestamp 1644511149
transform 1 0 26220 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_279
timestamp 1644511149
transform 1 0 26772 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_281
timestamp 1644511149
transform 1 0 26956 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_293
timestamp 1644511149
transform 1 0 28060 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_305
timestamp 1644511149
transform 1 0 29164 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_317
timestamp 1644511149
transform 1 0 30268 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_329
timestamp 1644511149
transform 1 0 31372 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_335
timestamp 1644511149
transform 1 0 31924 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_337
timestamp 1644511149
transform 1 0 32108 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_349
timestamp 1644511149
transform 1 0 33212 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_361
timestamp 1644511149
transform 1 0 34316 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_373
timestamp 1644511149
transform 1 0 35420 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_385
timestamp 1644511149
transform 1 0 36524 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_391
timestamp 1644511149
transform 1 0 37076 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_393
timestamp 1644511149
transform 1 0 37260 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_405
timestamp 1644511149
transform 1 0 38364 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_417
timestamp 1644511149
transform 1 0 39468 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_429
timestamp 1644511149
transform 1 0 40572 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_441
timestamp 1644511149
transform 1 0 41676 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_447
timestamp 1644511149
transform 1 0 42228 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_449
timestamp 1644511149
transform 1 0 42412 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_111_461
timestamp 1644511149
transform 1 0 43516 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_483
timestamp 1644511149
transform 1 0 45540 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_495
timestamp 1644511149
transform 1 0 46644 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_503
timestamp 1644511149
transform 1 0 47380 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_505
timestamp 1644511149
transform 1 0 47564 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_517
timestamp 1644511149
transform 1 0 48668 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_529
timestamp 1644511149
transform 1 0 49772 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_541
timestamp 1644511149
transform 1 0 50876 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_553
timestamp 1644511149
transform 1 0 51980 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_559
timestamp 1644511149
transform 1 0 52532 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_561
timestamp 1644511149
transform 1 0 52716 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_573
timestamp 1644511149
transform 1 0 53820 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_585
timestamp 1644511149
transform 1 0 54924 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_597
timestamp 1644511149
transform 1 0 56028 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_609
timestamp 1644511149
transform 1 0 57132 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_615
timestamp 1644511149
transform 1 0 57684 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_617
timestamp 1644511149
transform 1 0 57868 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_629
timestamp 1644511149
transform 1 0 58972 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_641
timestamp 1644511149
transform 1 0 60076 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_653
timestamp 1644511149
transform 1 0 61180 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_665
timestamp 1644511149
transform 1 0 62284 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_671
timestamp 1644511149
transform 1 0 62836 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_673
timestamp 1644511149
transform 1 0 63020 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_685
timestamp 1644511149
transform 1 0 64124 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_697
timestamp 1644511149
transform 1 0 65228 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_709
timestamp 1644511149
transform 1 0 66332 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_721
timestamp 1644511149
transform 1 0 67436 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_727
timestamp 1644511149
transform 1 0 67988 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_111_729
timestamp 1644511149
transform 1 0 68172 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_112_3
timestamp 1644511149
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_15
timestamp 1644511149
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1644511149
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_29
timestamp 1644511149
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_41
timestamp 1644511149
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_53
timestamp 1644511149
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_65
timestamp 1644511149
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1644511149
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1644511149
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_85
timestamp 1644511149
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_97
timestamp 1644511149
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_109
timestamp 1644511149
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_121
timestamp 1644511149
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_133
timestamp 1644511149
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_139
timestamp 1644511149
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_141
timestamp 1644511149
transform 1 0 14076 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_153
timestamp 1644511149
transform 1 0 15180 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_165
timestamp 1644511149
transform 1 0 16284 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_177
timestamp 1644511149
transform 1 0 17388 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_189
timestamp 1644511149
transform 1 0 18492 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_195
timestamp 1644511149
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_112_197
timestamp 1644511149
transform 1 0 19228 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_219
timestamp 1644511149
transform 1 0 21252 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_231
timestamp 1644511149
transform 1 0 22356 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_243
timestamp 1644511149
transform 1 0 23460 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_112_251
timestamp 1644511149
transform 1 0 24196 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_253
timestamp 1644511149
transform 1 0 24380 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_265
timestamp 1644511149
transform 1 0 25484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_277
timestamp 1644511149
transform 1 0 26588 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_289
timestamp 1644511149
transform 1 0 27692 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_301
timestamp 1644511149
transform 1 0 28796 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_307
timestamp 1644511149
transform 1 0 29348 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_309
timestamp 1644511149
transform 1 0 29532 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_321
timestamp 1644511149
transform 1 0 30636 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_333
timestamp 1644511149
transform 1 0 31740 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_345
timestamp 1644511149
transform 1 0 32844 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_357
timestamp 1644511149
transform 1 0 33948 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_363
timestamp 1644511149
transform 1 0 34500 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_365
timestamp 1644511149
transform 1 0 34684 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_377
timestamp 1644511149
transform 1 0 35788 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_389
timestamp 1644511149
transform 1 0 36892 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_401
timestamp 1644511149
transform 1 0 37996 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_413
timestamp 1644511149
transform 1 0 39100 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_419
timestamp 1644511149
transform 1 0 39652 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_421
timestamp 1644511149
transform 1 0 39836 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_433
timestamp 1644511149
transform 1 0 40940 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_445
timestamp 1644511149
transform 1 0 42044 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_112_457
timestamp 1644511149
transform 1 0 43148 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_112_462
timestamp 1644511149
transform 1 0 43608 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_112_469
timestamp 1644511149
transform 1 0 44252 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_475
timestamp 1644511149
transform 1 0 44804 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_477
timestamp 1644511149
transform 1 0 44988 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_489
timestamp 1644511149
transform 1 0 46092 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_501
timestamp 1644511149
transform 1 0 47196 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_513
timestamp 1644511149
transform 1 0 48300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_525
timestamp 1644511149
transform 1 0 49404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_531
timestamp 1644511149
transform 1 0 49956 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_533
timestamp 1644511149
transform 1 0 50140 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_545
timestamp 1644511149
transform 1 0 51244 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_557
timestamp 1644511149
transform 1 0 52348 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_569
timestamp 1644511149
transform 1 0 53452 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_581
timestamp 1644511149
transform 1 0 54556 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_587
timestamp 1644511149
transform 1 0 55108 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_589
timestamp 1644511149
transform 1 0 55292 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_601
timestamp 1644511149
transform 1 0 56396 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_613
timestamp 1644511149
transform 1 0 57500 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_625
timestamp 1644511149
transform 1 0 58604 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_637
timestamp 1644511149
transform 1 0 59708 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_643
timestamp 1644511149
transform 1 0 60260 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_645
timestamp 1644511149
transform 1 0 60444 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_657
timestamp 1644511149
transform 1 0 61548 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_669
timestamp 1644511149
transform 1 0 62652 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_681
timestamp 1644511149
transform 1 0 63756 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_693
timestamp 1644511149
transform 1 0 64860 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_699
timestamp 1644511149
transform 1 0 65412 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_701
timestamp 1644511149
transform 1 0 65596 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_713
timestamp 1644511149
transform 1 0 66700 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_725
timestamp 1644511149
transform 1 0 67804 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_3
timestamp 1644511149
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_15
timestamp 1644511149
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_27
timestamp 1644511149
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_39
timestamp 1644511149
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1644511149
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1644511149
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1644511149
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1644511149
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_81
timestamp 1644511149
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_93
timestamp 1644511149
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_105
timestamp 1644511149
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_111
timestamp 1644511149
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_113
timestamp 1644511149
transform 1 0 11500 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_125
timestamp 1644511149
transform 1 0 12604 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_137
timestamp 1644511149
transform 1 0 13708 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_149
timestamp 1644511149
transform 1 0 14812 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_161
timestamp 1644511149
transform 1 0 15916 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_167
timestamp 1644511149
transform 1 0 16468 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_169
timestamp 1644511149
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_181
timestamp 1644511149
transform 1 0 17756 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_113_189
timestamp 1644511149
transform 1 0 18492 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_113_195
timestamp 1644511149
transform 1 0 19044 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_220
timestamp 1644511149
transform 1 0 21344 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_113_225
timestamp 1644511149
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_237
timestamp 1644511149
transform 1 0 22908 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_249
timestamp 1644511149
transform 1 0 24012 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_261
timestamp 1644511149
transform 1 0 25116 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_273
timestamp 1644511149
transform 1 0 26220 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_279
timestamp 1644511149
transform 1 0 26772 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_281
timestamp 1644511149
transform 1 0 26956 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_293
timestamp 1644511149
transform 1 0 28060 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_305
timestamp 1644511149
transform 1 0 29164 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_317
timestamp 1644511149
transform 1 0 30268 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_329
timestamp 1644511149
transform 1 0 31372 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_335
timestamp 1644511149
transform 1 0 31924 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_337
timestamp 1644511149
transform 1 0 32108 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_349
timestamp 1644511149
transform 1 0 33212 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_361
timestamp 1644511149
transform 1 0 34316 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_373
timestamp 1644511149
transform 1 0 35420 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_385
timestamp 1644511149
transform 1 0 36524 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_391
timestamp 1644511149
transform 1 0 37076 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_393
timestamp 1644511149
transform 1 0 37260 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_405
timestamp 1644511149
transform 1 0 38364 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_417
timestamp 1644511149
transform 1 0 39468 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_429
timestamp 1644511149
transform 1 0 40572 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_441
timestamp 1644511149
transform 1 0 41676 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_447
timestamp 1644511149
transform 1 0 42228 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_449
timestamp 1644511149
transform 1 0 42412 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_461
timestamp 1644511149
transform 1 0 43516 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_473
timestamp 1644511149
transform 1 0 44620 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_485
timestamp 1644511149
transform 1 0 45724 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_497
timestamp 1644511149
transform 1 0 46828 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_503
timestamp 1644511149
transform 1 0 47380 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_505
timestamp 1644511149
transform 1 0 47564 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_517
timestamp 1644511149
transform 1 0 48668 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_529
timestamp 1644511149
transform 1 0 49772 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_541
timestamp 1644511149
transform 1 0 50876 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_553
timestamp 1644511149
transform 1 0 51980 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_559
timestamp 1644511149
transform 1 0 52532 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_561
timestamp 1644511149
transform 1 0 52716 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_573
timestamp 1644511149
transform 1 0 53820 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_585
timestamp 1644511149
transform 1 0 54924 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_597
timestamp 1644511149
transform 1 0 56028 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_609
timestamp 1644511149
transform 1 0 57132 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_615
timestamp 1644511149
transform 1 0 57684 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_617
timestamp 1644511149
transform 1 0 57868 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_629
timestamp 1644511149
transform 1 0 58972 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_641
timestamp 1644511149
transform 1 0 60076 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_653
timestamp 1644511149
transform 1 0 61180 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_665
timestamp 1644511149
transform 1 0 62284 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_671
timestamp 1644511149
transform 1 0 62836 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_673
timestamp 1644511149
transform 1 0 63020 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_685
timestamp 1644511149
transform 1 0 64124 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_697
timestamp 1644511149
transform 1 0 65228 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_709
timestamp 1644511149
transform 1 0 66332 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_721
timestamp 1644511149
transform 1 0 67436 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_727
timestamp 1644511149
transform 1 0 67988 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_113_729
timestamp 1644511149
transform 1 0 68172 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_114_3
timestamp 1644511149
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_15
timestamp 1644511149
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1644511149
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_29
timestamp 1644511149
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_41
timestamp 1644511149
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_53
timestamp 1644511149
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_65
timestamp 1644511149
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1644511149
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1644511149
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_85
timestamp 1644511149
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_97
timestamp 1644511149
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_109
timestamp 1644511149
transform 1 0 11132 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_121
timestamp 1644511149
transform 1 0 12236 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_133
timestamp 1644511149
transform 1 0 13340 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_139
timestamp 1644511149
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_141
timestamp 1644511149
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_153
timestamp 1644511149
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_165
timestamp 1644511149
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_177
timestamp 1644511149
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_189
timestamp 1644511149
transform 1 0 18492 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_195
timestamp 1644511149
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_114_197
timestamp 1644511149
transform 1 0 19228 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_114_206
timestamp 1644511149
transform 1 0 20056 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_218
timestamp 1644511149
transform 1 0 21160 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_230
timestamp 1644511149
transform 1 0 22264 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_242
timestamp 1644511149
transform 1 0 23368 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_114_250
timestamp 1644511149
transform 1 0 24104 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_114_253
timestamp 1644511149
transform 1 0 24380 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_265
timestamp 1644511149
transform 1 0 25484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_277
timestamp 1644511149
transform 1 0 26588 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_289
timestamp 1644511149
transform 1 0 27692 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_301
timestamp 1644511149
transform 1 0 28796 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_307
timestamp 1644511149
transform 1 0 29348 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_309
timestamp 1644511149
transform 1 0 29532 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_321
timestamp 1644511149
transform 1 0 30636 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_333
timestamp 1644511149
transform 1 0 31740 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_345
timestamp 1644511149
transform 1 0 32844 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_357
timestamp 1644511149
transform 1 0 33948 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_363
timestamp 1644511149
transform 1 0 34500 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_365
timestamp 1644511149
transform 1 0 34684 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_377
timestamp 1644511149
transform 1 0 35788 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_389
timestamp 1644511149
transform 1 0 36892 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_401
timestamp 1644511149
transform 1 0 37996 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_413
timestamp 1644511149
transform 1 0 39100 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_419
timestamp 1644511149
transform 1 0 39652 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_421
timestamp 1644511149
transform 1 0 39836 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_433
timestamp 1644511149
transform 1 0 40940 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_445
timestamp 1644511149
transform 1 0 42044 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_457
timestamp 1644511149
transform 1 0 43148 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_469
timestamp 1644511149
transform 1 0 44252 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_475
timestamp 1644511149
transform 1 0 44804 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_477
timestamp 1644511149
transform 1 0 44988 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_489
timestamp 1644511149
transform 1 0 46092 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_501
timestamp 1644511149
transform 1 0 47196 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_513
timestamp 1644511149
transform 1 0 48300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_525
timestamp 1644511149
transform 1 0 49404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_531
timestamp 1644511149
transform 1 0 49956 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_533
timestamp 1644511149
transform 1 0 50140 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_545
timestamp 1644511149
transform 1 0 51244 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_557
timestamp 1644511149
transform 1 0 52348 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_569
timestamp 1644511149
transform 1 0 53452 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_581
timestamp 1644511149
transform 1 0 54556 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_587
timestamp 1644511149
transform 1 0 55108 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_589
timestamp 1644511149
transform 1 0 55292 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_601
timestamp 1644511149
transform 1 0 56396 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_613
timestamp 1644511149
transform 1 0 57500 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_625
timestamp 1644511149
transform 1 0 58604 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_637
timestamp 1644511149
transform 1 0 59708 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_643
timestamp 1644511149
transform 1 0 60260 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_645
timestamp 1644511149
transform 1 0 60444 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_657
timestamp 1644511149
transform 1 0 61548 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_669
timestamp 1644511149
transform 1 0 62652 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_681
timestamp 1644511149
transform 1 0 63756 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_693
timestamp 1644511149
transform 1 0 64860 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_699
timestamp 1644511149
transform 1 0 65412 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_701
timestamp 1644511149
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_713
timestamp 1644511149
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_725
timestamp 1644511149
transform 1 0 67804 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_3
timestamp 1644511149
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_15
timestamp 1644511149
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_27
timestamp 1644511149
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_39
timestamp 1644511149
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1644511149
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1644511149
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_57
timestamp 1644511149
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_69
timestamp 1644511149
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_81
timestamp 1644511149
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_93
timestamp 1644511149
transform 1 0 9660 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_105
timestamp 1644511149
transform 1 0 10764 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_111
timestamp 1644511149
transform 1 0 11316 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_113
timestamp 1644511149
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_125
timestamp 1644511149
transform 1 0 12604 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_137
timestamp 1644511149
transform 1 0 13708 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_149
timestamp 1644511149
transform 1 0 14812 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_161
timestamp 1644511149
transform 1 0 15916 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_167
timestamp 1644511149
transform 1 0 16468 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_169
timestamp 1644511149
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_181
timestamp 1644511149
transform 1 0 17756 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_193
timestamp 1644511149
transform 1 0 18860 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_205
timestamp 1644511149
transform 1 0 19964 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_217
timestamp 1644511149
transform 1 0 21068 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_223
timestamp 1644511149
transform 1 0 21620 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_225
timestamp 1644511149
transform 1 0 21804 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_237
timestamp 1644511149
transform 1 0 22908 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_249
timestamp 1644511149
transform 1 0 24012 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_261
timestamp 1644511149
transform 1 0 25116 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_273
timestamp 1644511149
transform 1 0 26220 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_279
timestamp 1644511149
transform 1 0 26772 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_281
timestamp 1644511149
transform 1 0 26956 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_293
timestamp 1644511149
transform 1 0 28060 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_305
timestamp 1644511149
transform 1 0 29164 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_317
timestamp 1644511149
transform 1 0 30268 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_329
timestamp 1644511149
transform 1 0 31372 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_335
timestamp 1644511149
transform 1 0 31924 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_337
timestamp 1644511149
transform 1 0 32108 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_349
timestamp 1644511149
transform 1 0 33212 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_361
timestamp 1644511149
transform 1 0 34316 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_373
timestamp 1644511149
transform 1 0 35420 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_385
timestamp 1644511149
transform 1 0 36524 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_391
timestamp 1644511149
transform 1 0 37076 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_393
timestamp 1644511149
transform 1 0 37260 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_405
timestamp 1644511149
transform 1 0 38364 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_417
timestamp 1644511149
transform 1 0 39468 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_429
timestamp 1644511149
transform 1 0 40572 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_441
timestamp 1644511149
transform 1 0 41676 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_447
timestamp 1644511149
transform 1 0 42228 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_449
timestamp 1644511149
transform 1 0 42412 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_461
timestamp 1644511149
transform 1 0 43516 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_473
timestamp 1644511149
transform 1 0 44620 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_485
timestamp 1644511149
transform 1 0 45724 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_497
timestamp 1644511149
transform 1 0 46828 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_503
timestamp 1644511149
transform 1 0 47380 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_505
timestamp 1644511149
transform 1 0 47564 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_517
timestamp 1644511149
transform 1 0 48668 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_529
timestamp 1644511149
transform 1 0 49772 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_541
timestamp 1644511149
transform 1 0 50876 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_553
timestamp 1644511149
transform 1 0 51980 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_559
timestamp 1644511149
transform 1 0 52532 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_561
timestamp 1644511149
transform 1 0 52716 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_573
timestamp 1644511149
transform 1 0 53820 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_585
timestamp 1644511149
transform 1 0 54924 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_597
timestamp 1644511149
transform 1 0 56028 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_609
timestamp 1644511149
transform 1 0 57132 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_615
timestamp 1644511149
transform 1 0 57684 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_617
timestamp 1644511149
transform 1 0 57868 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_629
timestamp 1644511149
transform 1 0 58972 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_641
timestamp 1644511149
transform 1 0 60076 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_653
timestamp 1644511149
transform 1 0 61180 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_665
timestamp 1644511149
transform 1 0 62284 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_671
timestamp 1644511149
transform 1 0 62836 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_673
timestamp 1644511149
transform 1 0 63020 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_685
timestamp 1644511149
transform 1 0 64124 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_697
timestamp 1644511149
transform 1 0 65228 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_709
timestamp 1644511149
transform 1 0 66332 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_721
timestamp 1644511149
transform 1 0 67436 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_727
timestamp 1644511149
transform 1 0 67988 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_115_729
timestamp 1644511149
transform 1 0 68172 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_3
timestamp 1644511149
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_15
timestamp 1644511149
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1644511149
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_29
timestamp 1644511149
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_41
timestamp 1644511149
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_53
timestamp 1644511149
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_65
timestamp 1644511149
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_77
timestamp 1644511149
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1644511149
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_85
timestamp 1644511149
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_97
timestamp 1644511149
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_109
timestamp 1644511149
transform 1 0 11132 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_121
timestamp 1644511149
transform 1 0 12236 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_133
timestamp 1644511149
transform 1 0 13340 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_139
timestamp 1644511149
transform 1 0 13892 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_141
timestamp 1644511149
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_153
timestamp 1644511149
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_165
timestamp 1644511149
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_177
timestamp 1644511149
transform 1 0 17388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_189
timestamp 1644511149
transform 1 0 18492 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_195
timestamp 1644511149
transform 1 0 19044 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_197
timestamp 1644511149
transform 1 0 19228 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_209
timestamp 1644511149
transform 1 0 20332 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_221
timestamp 1644511149
transform 1 0 21436 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_233
timestamp 1644511149
transform 1 0 22540 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_245
timestamp 1644511149
transform 1 0 23644 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_251
timestamp 1644511149
transform 1 0 24196 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_253
timestamp 1644511149
transform 1 0 24380 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_265
timestamp 1644511149
transform 1 0 25484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_277
timestamp 1644511149
transform 1 0 26588 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_289
timestamp 1644511149
transform 1 0 27692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_301
timestamp 1644511149
transform 1 0 28796 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_307
timestamp 1644511149
transform 1 0 29348 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_309
timestamp 1644511149
transform 1 0 29532 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_321
timestamp 1644511149
transform 1 0 30636 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_333
timestamp 1644511149
transform 1 0 31740 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_345
timestamp 1644511149
transform 1 0 32844 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_357
timestamp 1644511149
transform 1 0 33948 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_363
timestamp 1644511149
transform 1 0 34500 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_365
timestamp 1644511149
transform 1 0 34684 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_377
timestamp 1644511149
transform 1 0 35788 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_389
timestamp 1644511149
transform 1 0 36892 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_401
timestamp 1644511149
transform 1 0 37996 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_413
timestamp 1644511149
transform 1 0 39100 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_419
timestamp 1644511149
transform 1 0 39652 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_421
timestamp 1644511149
transform 1 0 39836 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_433
timestamp 1644511149
transform 1 0 40940 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_445
timestamp 1644511149
transform 1 0 42044 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_457
timestamp 1644511149
transform 1 0 43148 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_469
timestamp 1644511149
transform 1 0 44252 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_475
timestamp 1644511149
transform 1 0 44804 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_477
timestamp 1644511149
transform 1 0 44988 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_489
timestamp 1644511149
transform 1 0 46092 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_501
timestamp 1644511149
transform 1 0 47196 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_513
timestamp 1644511149
transform 1 0 48300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_525
timestamp 1644511149
transform 1 0 49404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_531
timestamp 1644511149
transform 1 0 49956 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_533
timestamp 1644511149
transform 1 0 50140 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_545
timestamp 1644511149
transform 1 0 51244 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_557
timestamp 1644511149
transform 1 0 52348 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_569
timestamp 1644511149
transform 1 0 53452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_581
timestamp 1644511149
transform 1 0 54556 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_587
timestamp 1644511149
transform 1 0 55108 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_589
timestamp 1644511149
transform 1 0 55292 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_601
timestamp 1644511149
transform 1 0 56396 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_613
timestamp 1644511149
transform 1 0 57500 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_625
timestamp 1644511149
transform 1 0 58604 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_637
timestamp 1644511149
transform 1 0 59708 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_643
timestamp 1644511149
transform 1 0 60260 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_645
timestamp 1644511149
transform 1 0 60444 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_657
timestamp 1644511149
transform 1 0 61548 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_669
timestamp 1644511149
transform 1 0 62652 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_681
timestamp 1644511149
transform 1 0 63756 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_693
timestamp 1644511149
transform 1 0 64860 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_699
timestamp 1644511149
transform 1 0 65412 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_701
timestamp 1644511149
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_713
timestamp 1644511149
transform 1 0 66700 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_725
timestamp 1644511149
transform 1 0 67804 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_9
timestamp 1644511149
transform 1 0 1932 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_21
timestamp 1644511149
transform 1 0 3036 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_33
timestamp 1644511149
transform 1 0 4140 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_45
timestamp 1644511149
transform 1 0 5244 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_117_53
timestamp 1644511149
transform 1 0 5980 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1644511149
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1644511149
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_81
timestamp 1644511149
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_93
timestamp 1644511149
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_105
timestamp 1644511149
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_111
timestamp 1644511149
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_113
timestamp 1644511149
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_125
timestamp 1644511149
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_137
timestamp 1644511149
transform 1 0 13708 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_149
timestamp 1644511149
transform 1 0 14812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_161
timestamp 1644511149
transform 1 0 15916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_167
timestamp 1644511149
transform 1 0 16468 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_169
timestamp 1644511149
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_181
timestamp 1644511149
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_193
timestamp 1644511149
transform 1 0 18860 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_205
timestamp 1644511149
transform 1 0 19964 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_217
timestamp 1644511149
transform 1 0 21068 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_223
timestamp 1644511149
transform 1 0 21620 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_225
timestamp 1644511149
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_237
timestamp 1644511149
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_249
timestamp 1644511149
transform 1 0 24012 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_261
timestamp 1644511149
transform 1 0 25116 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_273
timestamp 1644511149
transform 1 0 26220 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_279
timestamp 1644511149
transform 1 0 26772 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_281
timestamp 1644511149
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_293
timestamp 1644511149
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_305
timestamp 1644511149
transform 1 0 29164 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_317
timestamp 1644511149
transform 1 0 30268 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_329
timestamp 1644511149
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_335
timestamp 1644511149
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_337
timestamp 1644511149
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_349
timestamp 1644511149
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_361
timestamp 1644511149
transform 1 0 34316 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_373
timestamp 1644511149
transform 1 0 35420 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_385
timestamp 1644511149
transform 1 0 36524 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_391
timestamp 1644511149
transform 1 0 37076 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_393
timestamp 1644511149
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_405
timestamp 1644511149
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_417
timestamp 1644511149
transform 1 0 39468 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_429
timestamp 1644511149
transform 1 0 40572 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_441
timestamp 1644511149
transform 1 0 41676 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_447
timestamp 1644511149
transform 1 0 42228 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_449
timestamp 1644511149
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_461
timestamp 1644511149
transform 1 0 43516 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_473
timestamp 1644511149
transform 1 0 44620 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_485
timestamp 1644511149
transform 1 0 45724 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_497
timestamp 1644511149
transform 1 0 46828 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_503
timestamp 1644511149
transform 1 0 47380 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_505
timestamp 1644511149
transform 1 0 47564 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_517
timestamp 1644511149
transform 1 0 48668 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_529
timestamp 1644511149
transform 1 0 49772 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_541
timestamp 1644511149
transform 1 0 50876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_553
timestamp 1644511149
transform 1 0 51980 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_559
timestamp 1644511149
transform 1 0 52532 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_561
timestamp 1644511149
transform 1 0 52716 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_573
timestamp 1644511149
transform 1 0 53820 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_585
timestamp 1644511149
transform 1 0 54924 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_597
timestamp 1644511149
transform 1 0 56028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_609
timestamp 1644511149
transform 1 0 57132 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_615
timestamp 1644511149
transform 1 0 57684 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_617
timestamp 1644511149
transform 1 0 57868 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_629
timestamp 1644511149
transform 1 0 58972 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_641
timestamp 1644511149
transform 1 0 60076 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_653
timestamp 1644511149
transform 1 0 61180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_665
timestamp 1644511149
transform 1 0 62284 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_671
timestamp 1644511149
transform 1 0 62836 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_673
timestamp 1644511149
transform 1 0 63020 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_685
timestamp 1644511149
transform 1 0 64124 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_697
timestamp 1644511149
transform 1 0 65228 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_709
timestamp 1644511149
transform 1 0 66332 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_721
timestamp 1644511149
transform 1 0 67436 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_727
timestamp 1644511149
transform 1 0 67988 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_729
timestamp 1644511149
transform 1 0 68172 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_118_3
timestamp 1644511149
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_15
timestamp 1644511149
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1644511149
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_29
timestamp 1644511149
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_41
timestamp 1644511149
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_53
timestamp 1644511149
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_65
timestamp 1644511149
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1644511149
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1644511149
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_85
timestamp 1644511149
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_97
timestamp 1644511149
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_109
timestamp 1644511149
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_121
timestamp 1644511149
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1644511149
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1644511149
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_141
timestamp 1644511149
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_153
timestamp 1644511149
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_165
timestamp 1644511149
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_177
timestamp 1644511149
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1644511149
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1644511149
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_197
timestamp 1644511149
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_209
timestamp 1644511149
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_221
timestamp 1644511149
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_233
timestamp 1644511149
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_245
timestamp 1644511149
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1644511149
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_253
timestamp 1644511149
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_265
timestamp 1644511149
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_277
timestamp 1644511149
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_289
timestamp 1644511149
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_301
timestamp 1644511149
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_307
timestamp 1644511149
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_309
timestamp 1644511149
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_321
timestamp 1644511149
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_333
timestamp 1644511149
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_345
timestamp 1644511149
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_357
timestamp 1644511149
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_363
timestamp 1644511149
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_365
timestamp 1644511149
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_377
timestamp 1644511149
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_389
timestamp 1644511149
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_401
timestamp 1644511149
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_413
timestamp 1644511149
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1644511149
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_421
timestamp 1644511149
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_433
timestamp 1644511149
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_445
timestamp 1644511149
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_457
timestamp 1644511149
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_469
timestamp 1644511149
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_475
timestamp 1644511149
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_477
timestamp 1644511149
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_489
timestamp 1644511149
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_501
timestamp 1644511149
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_513
timestamp 1644511149
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_525
timestamp 1644511149
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_531
timestamp 1644511149
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_533
timestamp 1644511149
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_545
timestamp 1644511149
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_557
timestamp 1644511149
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_569
timestamp 1644511149
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_581
timestamp 1644511149
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1644511149
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_589
timestamp 1644511149
transform 1 0 55292 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_601
timestamp 1644511149
transform 1 0 56396 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_613
timestamp 1644511149
transform 1 0 57500 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_625
timestamp 1644511149
transform 1 0 58604 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_637
timestamp 1644511149
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_643
timestamp 1644511149
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_645
timestamp 1644511149
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_657
timestamp 1644511149
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_669
timestamp 1644511149
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_681
timestamp 1644511149
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_693
timestamp 1644511149
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1644511149
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_701
timestamp 1644511149
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_713
timestamp 1644511149
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_725
timestamp 1644511149
transform 1 0 67804 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_3
timestamp 1644511149
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_15
timestamp 1644511149
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_27
timestamp 1644511149
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_39
timestamp 1644511149
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1644511149
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1644511149
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1644511149
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_69
timestamp 1644511149
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_81
timestamp 1644511149
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_93
timestamp 1644511149
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1644511149
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1644511149
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_113
timestamp 1644511149
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_125
timestamp 1644511149
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_137
timestamp 1644511149
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_149
timestamp 1644511149
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1644511149
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1644511149
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_169
timestamp 1644511149
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_181
timestamp 1644511149
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_193
timestamp 1644511149
transform 1 0 18860 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_205
timestamp 1644511149
transform 1 0 19964 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_217
timestamp 1644511149
transform 1 0 21068 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1644511149
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_225
timestamp 1644511149
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_237
timestamp 1644511149
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_249
timestamp 1644511149
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_261
timestamp 1644511149
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_273
timestamp 1644511149
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1644511149
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_281
timestamp 1644511149
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_293
timestamp 1644511149
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_305
timestamp 1644511149
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_317
timestamp 1644511149
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_329
timestamp 1644511149
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_335
timestamp 1644511149
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_337
timestamp 1644511149
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_349
timestamp 1644511149
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_361
timestamp 1644511149
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_373
timestamp 1644511149
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_385
timestamp 1644511149
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_391
timestamp 1644511149
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_393
timestamp 1644511149
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_405
timestamp 1644511149
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_417
timestamp 1644511149
transform 1 0 39468 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_429
timestamp 1644511149
transform 1 0 40572 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_441
timestamp 1644511149
transform 1 0 41676 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_447
timestamp 1644511149
transform 1 0 42228 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_449
timestamp 1644511149
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_461
timestamp 1644511149
transform 1 0 43516 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_473
timestamp 1644511149
transform 1 0 44620 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_485
timestamp 1644511149
transform 1 0 45724 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_497
timestamp 1644511149
transform 1 0 46828 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1644511149
transform 1 0 47380 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_505
timestamp 1644511149
transform 1 0 47564 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_517
timestamp 1644511149
transform 1 0 48668 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_529
timestamp 1644511149
transform 1 0 49772 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_541
timestamp 1644511149
transform 1 0 50876 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_553
timestamp 1644511149
transform 1 0 51980 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_559
timestamp 1644511149
transform 1 0 52532 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_561
timestamp 1644511149
transform 1 0 52716 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_573
timestamp 1644511149
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_585
timestamp 1644511149
transform 1 0 54924 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_597
timestamp 1644511149
transform 1 0 56028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_609
timestamp 1644511149
transform 1 0 57132 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_615
timestamp 1644511149
transform 1 0 57684 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_617
timestamp 1644511149
transform 1 0 57868 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_629
timestamp 1644511149
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_641
timestamp 1644511149
transform 1 0 60076 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_653
timestamp 1644511149
transform 1 0 61180 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_665
timestamp 1644511149
transform 1 0 62284 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_671
timestamp 1644511149
transform 1 0 62836 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_673
timestamp 1644511149
transform 1 0 63020 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_685
timestamp 1644511149
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_697
timestamp 1644511149
transform 1 0 65228 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_709
timestamp 1644511149
transform 1 0 66332 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_721
timestamp 1644511149
transform 1 0 67436 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_727
timestamp 1644511149
transform 1 0 67988 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_729
timestamp 1644511149
transform 1 0 68172 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_120_3
timestamp 1644511149
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_15
timestamp 1644511149
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1644511149
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_29
timestamp 1644511149
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_41
timestamp 1644511149
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_53
timestamp 1644511149
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_65
timestamp 1644511149
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1644511149
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1644511149
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_85
timestamp 1644511149
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_97
timestamp 1644511149
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_109
timestamp 1644511149
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_121
timestamp 1644511149
transform 1 0 12236 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_133
timestamp 1644511149
transform 1 0 13340 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1644511149
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_141
timestamp 1644511149
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_153
timestamp 1644511149
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_165
timestamp 1644511149
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_177
timestamp 1644511149
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_189
timestamp 1644511149
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_195
timestamp 1644511149
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_197
timestamp 1644511149
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_209
timestamp 1644511149
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_221
timestamp 1644511149
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_233
timestamp 1644511149
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1644511149
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1644511149
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_253
timestamp 1644511149
transform 1 0 24380 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_265
timestamp 1644511149
transform 1 0 25484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_277
timestamp 1644511149
transform 1 0 26588 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_289
timestamp 1644511149
transform 1 0 27692 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_301
timestamp 1644511149
transform 1 0 28796 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_307
timestamp 1644511149
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_309
timestamp 1644511149
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_321
timestamp 1644511149
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_333
timestamp 1644511149
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_345
timestamp 1644511149
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_357
timestamp 1644511149
transform 1 0 33948 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1644511149
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_365
timestamp 1644511149
transform 1 0 34684 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_377
timestamp 1644511149
transform 1 0 35788 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_389
timestamp 1644511149
transform 1 0 36892 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_401
timestamp 1644511149
transform 1 0 37996 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_413
timestamp 1644511149
transform 1 0 39100 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_419
timestamp 1644511149
transform 1 0 39652 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_421
timestamp 1644511149
transform 1 0 39836 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_433
timestamp 1644511149
transform 1 0 40940 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_445
timestamp 1644511149
transform 1 0 42044 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_457
timestamp 1644511149
transform 1 0 43148 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_469
timestamp 1644511149
transform 1 0 44252 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_475
timestamp 1644511149
transform 1 0 44804 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_477
timestamp 1644511149
transform 1 0 44988 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_489
timestamp 1644511149
transform 1 0 46092 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_501
timestamp 1644511149
transform 1 0 47196 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_513
timestamp 1644511149
transform 1 0 48300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_525
timestamp 1644511149
transform 1 0 49404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_531
timestamp 1644511149
transform 1 0 49956 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_533
timestamp 1644511149
transform 1 0 50140 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_545
timestamp 1644511149
transform 1 0 51244 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_557
timestamp 1644511149
transform 1 0 52348 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_569
timestamp 1644511149
transform 1 0 53452 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_581
timestamp 1644511149
transform 1 0 54556 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_587
timestamp 1644511149
transform 1 0 55108 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_589
timestamp 1644511149
transform 1 0 55292 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_601
timestamp 1644511149
transform 1 0 56396 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_613
timestamp 1644511149
transform 1 0 57500 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_625
timestamp 1644511149
transform 1 0 58604 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_637
timestamp 1644511149
transform 1 0 59708 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_643
timestamp 1644511149
transform 1 0 60260 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_645
timestamp 1644511149
transform 1 0 60444 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_657
timestamp 1644511149
transform 1 0 61548 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_669
timestamp 1644511149
transform 1 0 62652 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_681
timestamp 1644511149
transform 1 0 63756 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_693
timestamp 1644511149
transform 1 0 64860 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_699
timestamp 1644511149
transform 1 0 65412 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_701
timestamp 1644511149
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_713
timestamp 1644511149
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_725
timestamp 1644511149
transform 1 0 67804 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_121_3
timestamp 1644511149
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_15
timestamp 1644511149
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_27
timestamp 1644511149
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_39
timestamp 1644511149
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1644511149
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1644511149
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1644511149
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1644511149
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_81
timestamp 1644511149
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_93
timestamp 1644511149
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1644511149
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1644511149
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_113
timestamp 1644511149
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_125
timestamp 1644511149
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_137
timestamp 1644511149
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_149
timestamp 1644511149
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1644511149
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1644511149
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_169
timestamp 1644511149
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_181
timestamp 1644511149
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_193
timestamp 1644511149
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_205
timestamp 1644511149
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_217
timestamp 1644511149
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_223
timestamp 1644511149
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_225
timestamp 1644511149
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_237
timestamp 1644511149
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_249
timestamp 1644511149
transform 1 0 24012 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_261
timestamp 1644511149
transform 1 0 25116 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_273
timestamp 1644511149
transform 1 0 26220 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1644511149
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_281
timestamp 1644511149
transform 1 0 26956 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_293
timestamp 1644511149
transform 1 0 28060 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_305
timestamp 1644511149
transform 1 0 29164 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_317
timestamp 1644511149
transform 1 0 30268 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_329
timestamp 1644511149
transform 1 0 31372 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_335
timestamp 1644511149
transform 1 0 31924 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_337
timestamp 1644511149
transform 1 0 32108 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_349
timestamp 1644511149
transform 1 0 33212 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_361
timestamp 1644511149
transform 1 0 34316 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_373
timestamp 1644511149
transform 1 0 35420 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_385
timestamp 1644511149
transform 1 0 36524 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_391
timestamp 1644511149
transform 1 0 37076 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_393
timestamp 1644511149
transform 1 0 37260 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_405
timestamp 1644511149
transform 1 0 38364 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_417
timestamp 1644511149
transform 1 0 39468 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_429
timestamp 1644511149
transform 1 0 40572 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_441
timestamp 1644511149
transform 1 0 41676 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_447
timestamp 1644511149
transform 1 0 42228 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_449
timestamp 1644511149
transform 1 0 42412 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_461
timestamp 1644511149
transform 1 0 43516 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_473
timestamp 1644511149
transform 1 0 44620 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_485
timestamp 1644511149
transform 1 0 45724 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_497
timestamp 1644511149
transform 1 0 46828 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_503
timestamp 1644511149
transform 1 0 47380 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_505
timestamp 1644511149
transform 1 0 47564 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_517
timestamp 1644511149
transform 1 0 48668 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_529
timestamp 1644511149
transform 1 0 49772 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_541
timestamp 1644511149
transform 1 0 50876 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_553
timestamp 1644511149
transform 1 0 51980 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_559
timestamp 1644511149
transform 1 0 52532 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_561
timestamp 1644511149
transform 1 0 52716 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_573
timestamp 1644511149
transform 1 0 53820 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_585
timestamp 1644511149
transform 1 0 54924 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_597
timestamp 1644511149
transform 1 0 56028 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_609
timestamp 1644511149
transform 1 0 57132 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_615
timestamp 1644511149
transform 1 0 57684 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_617
timestamp 1644511149
transform 1 0 57868 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_629
timestamp 1644511149
transform 1 0 58972 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_641
timestamp 1644511149
transform 1 0 60076 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_653
timestamp 1644511149
transform 1 0 61180 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_665
timestamp 1644511149
transform 1 0 62284 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_671
timestamp 1644511149
transform 1 0 62836 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_673
timestamp 1644511149
transform 1 0 63020 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_685
timestamp 1644511149
transform 1 0 64124 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_697
timestamp 1644511149
transform 1 0 65228 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_709
timestamp 1644511149
transform 1 0 66332 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_721
timestamp 1644511149
transform 1 0 67436 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_727
timestamp 1644511149
transform 1 0 67988 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_121_729
timestamp 1644511149
transform 1 0 68172 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_122_3
timestamp 1644511149
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_15
timestamp 1644511149
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1644511149
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_29
timestamp 1644511149
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_41
timestamp 1644511149
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_53
timestamp 1644511149
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_65
timestamp 1644511149
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1644511149
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1644511149
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_85
timestamp 1644511149
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_97
timestamp 1644511149
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_109
timestamp 1644511149
transform 1 0 11132 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_121
timestamp 1644511149
transform 1 0 12236 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_133
timestamp 1644511149
transform 1 0 13340 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_139
timestamp 1644511149
transform 1 0 13892 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_141
timestamp 1644511149
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_153
timestamp 1644511149
transform 1 0 15180 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_165
timestamp 1644511149
transform 1 0 16284 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_177
timestamp 1644511149
transform 1 0 17388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_189
timestamp 1644511149
transform 1 0 18492 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_195
timestamp 1644511149
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_197
timestamp 1644511149
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_209
timestamp 1644511149
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_221
timestamp 1644511149
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_233
timestamp 1644511149
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_245
timestamp 1644511149
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_251
timestamp 1644511149
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_253
timestamp 1644511149
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_265
timestamp 1644511149
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_277
timestamp 1644511149
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_289
timestamp 1644511149
transform 1 0 27692 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_301
timestamp 1644511149
transform 1 0 28796 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_307
timestamp 1644511149
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_309
timestamp 1644511149
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_321
timestamp 1644511149
transform 1 0 30636 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_333
timestamp 1644511149
transform 1 0 31740 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_345
timestamp 1644511149
transform 1 0 32844 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_357
timestamp 1644511149
transform 1 0 33948 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_363
timestamp 1644511149
transform 1 0 34500 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_365
timestamp 1644511149
transform 1 0 34684 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_377
timestamp 1644511149
transform 1 0 35788 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_389
timestamp 1644511149
transform 1 0 36892 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_401
timestamp 1644511149
transform 1 0 37996 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_413
timestamp 1644511149
transform 1 0 39100 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_419
timestamp 1644511149
transform 1 0 39652 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_421
timestamp 1644511149
transform 1 0 39836 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_433
timestamp 1644511149
transform 1 0 40940 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_445
timestamp 1644511149
transform 1 0 42044 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_457
timestamp 1644511149
transform 1 0 43148 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_469
timestamp 1644511149
transform 1 0 44252 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_475
timestamp 1644511149
transform 1 0 44804 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_477
timestamp 1644511149
transform 1 0 44988 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_489
timestamp 1644511149
transform 1 0 46092 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_501
timestamp 1644511149
transform 1 0 47196 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_513
timestamp 1644511149
transform 1 0 48300 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_525
timestamp 1644511149
transform 1 0 49404 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_531
timestamp 1644511149
transform 1 0 49956 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_533
timestamp 1644511149
transform 1 0 50140 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_545
timestamp 1644511149
transform 1 0 51244 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_557
timestamp 1644511149
transform 1 0 52348 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_569
timestamp 1644511149
transform 1 0 53452 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_581
timestamp 1644511149
transform 1 0 54556 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_587
timestamp 1644511149
transform 1 0 55108 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_589
timestamp 1644511149
transform 1 0 55292 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_601
timestamp 1644511149
transform 1 0 56396 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_613
timestamp 1644511149
transform 1 0 57500 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_625
timestamp 1644511149
transform 1 0 58604 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_637
timestamp 1644511149
transform 1 0 59708 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_643
timestamp 1644511149
transform 1 0 60260 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_645
timestamp 1644511149
transform 1 0 60444 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_657
timestamp 1644511149
transform 1 0 61548 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_669
timestamp 1644511149
transform 1 0 62652 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_681
timestamp 1644511149
transform 1 0 63756 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_693
timestamp 1644511149
transform 1 0 64860 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_699
timestamp 1644511149
transform 1 0 65412 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_701
timestamp 1644511149
transform 1 0 65596 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_713
timestamp 1644511149
transform 1 0 66700 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_725
timestamp 1644511149
transform 1 0 67804 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_123_3
timestamp 1644511149
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_15
timestamp 1644511149
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_123_27
timestamp 1644511149
transform 1 0 3588 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_29
timestamp 1644511149
transform 1 0 3772 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_41
timestamp 1644511149
transform 1 0 4876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_53
timestamp 1644511149
transform 1 0 5980 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_57
timestamp 1644511149
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_69
timestamp 1644511149
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_81
timestamp 1644511149
transform 1 0 8556 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_85
timestamp 1644511149
transform 1 0 8924 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_97
timestamp 1644511149
transform 1 0 10028 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_109
timestamp 1644511149
transform 1 0 11132 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_113
timestamp 1644511149
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_125
timestamp 1644511149
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_137
timestamp 1644511149
transform 1 0 13708 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_141
timestamp 1644511149
transform 1 0 14076 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_153
timestamp 1644511149
transform 1 0 15180 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_165
timestamp 1644511149
transform 1 0 16284 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_169
timestamp 1644511149
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_181
timestamp 1644511149
transform 1 0 17756 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_193
timestamp 1644511149
transform 1 0 18860 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_197
timestamp 1644511149
transform 1 0 19228 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_209
timestamp 1644511149
transform 1 0 20332 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_221
timestamp 1644511149
transform 1 0 21436 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_225
timestamp 1644511149
transform 1 0 21804 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_237
timestamp 1644511149
transform 1 0 22908 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_249
timestamp 1644511149
transform 1 0 24012 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_253
timestamp 1644511149
transform 1 0 24380 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_265
timestamp 1644511149
transform 1 0 25484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_277
timestamp 1644511149
transform 1 0 26588 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_281
timestamp 1644511149
transform 1 0 26956 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_293
timestamp 1644511149
transform 1 0 28060 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_305
timestamp 1644511149
transform 1 0 29164 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_309
timestamp 1644511149
transform 1 0 29532 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_321
timestamp 1644511149
transform 1 0 30636 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_333
timestamp 1644511149
transform 1 0 31740 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_337
timestamp 1644511149
transform 1 0 32108 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_349
timestamp 1644511149
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_361
timestamp 1644511149
transform 1 0 34316 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_365
timestamp 1644511149
transform 1 0 34684 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_377
timestamp 1644511149
transform 1 0 35788 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_389
timestamp 1644511149
transform 1 0 36892 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_393
timestamp 1644511149
transform 1 0 37260 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_405
timestamp 1644511149
transform 1 0 38364 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_417
timestamp 1644511149
transform 1 0 39468 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_421
timestamp 1644511149
transform 1 0 39836 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_433
timestamp 1644511149
transform 1 0 40940 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_445
timestamp 1644511149
transform 1 0 42044 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_449
timestamp 1644511149
transform 1 0 42412 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_461
timestamp 1644511149
transform 1 0 43516 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_473
timestamp 1644511149
transform 1 0 44620 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_477
timestamp 1644511149
transform 1 0 44988 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_489
timestamp 1644511149
transform 1 0 46092 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_501
timestamp 1644511149
transform 1 0 47196 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_505
timestamp 1644511149
transform 1 0 47564 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_517
timestamp 1644511149
transform 1 0 48668 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_529
timestamp 1644511149
transform 1 0 49772 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_533
timestamp 1644511149
transform 1 0 50140 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_545
timestamp 1644511149
transform 1 0 51244 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_557
timestamp 1644511149
transform 1 0 52348 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_561
timestamp 1644511149
transform 1 0 52716 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_573
timestamp 1644511149
transform 1 0 53820 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_585
timestamp 1644511149
transform 1 0 54924 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_589
timestamp 1644511149
transform 1 0 55292 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_601
timestamp 1644511149
transform 1 0 56396 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_613
timestamp 1644511149
transform 1 0 57500 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_617
timestamp 1644511149
transform 1 0 57868 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_629
timestamp 1644511149
transform 1 0 58972 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_641
timestamp 1644511149
transform 1 0 60076 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_645
timestamp 1644511149
transform 1 0 60444 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_657
timestamp 1644511149
transform 1 0 61548 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_669
timestamp 1644511149
transform 1 0 62652 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_673
timestamp 1644511149
transform 1 0 63020 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_685
timestamp 1644511149
transform 1 0 64124 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_697
timestamp 1644511149
transform 1 0 65228 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_701
timestamp 1644511149
transform 1 0 65596 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_713
timestamp 1644511149
transform 1 0 66700 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_725
timestamp 1644511149
transform 1 0 67804 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_123_729
timestamp 1644511149
transform 1 0 68172 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 68816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 68816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 68816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 68816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 68816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 68816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 68816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 68816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 68816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 68816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 68816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 68816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 68816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 68816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 68816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 68816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 68816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 68816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 68816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 68816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 68816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 68816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 68816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 68816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 68816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 68816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 68816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 68816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 68816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 68816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 68816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 68816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 68816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 68816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 68816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 68816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 68816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 68816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 68816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 68816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 68816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 68816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 68816 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 68816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 68816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 68816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 68816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 68816 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 68816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 68816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 68816 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 68816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 68816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 68816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 68816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 68816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 68816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 68816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 68816 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 68816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 68816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 68816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 68816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 68816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 68816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 68816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 68816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 68816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 68816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 68816 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 68816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 68816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 68816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 68816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 68816 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 68816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 68816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 68816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 68816 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 68816 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1644511149
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1644511149
transform -1 0 68816 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1644511149
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1644511149
transform -1 0 68816 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1644511149
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1644511149
transform -1 0 68816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1644511149
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1644511149
transform -1 0 68816 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1644511149
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1644511149
transform -1 0 68816 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1644511149
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1644511149
transform -1 0 68816 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1644511149
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1644511149
transform -1 0 68816 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1644511149
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1644511149
transform -1 0 68816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1644511149
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1644511149
transform -1 0 68816 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1644511149
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1644511149
transform -1 0 68816 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1644511149
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1644511149
transform -1 0 68816 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1644511149
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1644511149
transform -1 0 68816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1644511149
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1644511149
transform -1 0 68816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1644511149
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1644511149
transform -1 0 68816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1644511149
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1644511149
transform -1 0 68816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1644511149
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1644511149
transform -1 0 68816 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1644511149
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1644511149
transform -1 0 68816 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1644511149
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1644511149
transform -1 0 68816 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1644511149
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1644511149
transform -1 0 68816 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1644511149
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1644511149
transform -1 0 68816 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1644511149
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1644511149
transform -1 0 68816 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1644511149
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1644511149
transform -1 0 68816 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1644511149
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1644511149
transform -1 0 68816 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1644511149
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1644511149
transform -1 0 68816 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1644511149
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1644511149
transform -1 0 68816 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1644511149
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1644511149
transform -1 0 68816 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1644511149
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1644511149
transform -1 0 68816 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1644511149
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1644511149
transform -1 0 68816 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1644511149
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1644511149
transform -1 0 68816 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1644511149
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1644511149
transform -1 0 68816 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1644511149
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1644511149
transform -1 0 68816 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1644511149
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1644511149
transform -1 0 68816 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1644511149
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1644511149
transform -1 0 68816 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1644511149
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1644511149
transform -1 0 68816 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1644511149
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1644511149
transform -1 0 68816 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1644511149
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1644511149
transform -1 0 68816 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1644511149
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1644511149
transform -1 0 68816 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1644511149
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1644511149
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1644511149
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1644511149
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1644511149
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1644511149
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1644511149
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1644511149
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1644511149
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1644511149
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1644511149
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1644511149
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1644511149
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1644511149
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1644511149
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1644511149
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1644511149
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1644511149
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1644511149
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1644511149
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1644511149
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1644511149
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1644511149
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1644511149
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1644511149
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1644511149
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1644511149
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1644511149
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1644511149
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1644511149
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1644511149
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1644511149
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1644511149
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1644511149
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1644511149
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1644511149
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1644511149
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1644511149
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1644511149
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1644511149
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1644511149
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1644511149
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1644511149
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1644511149
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1644511149
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1644511149
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1644511149
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1644511149
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1644511149
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1644511149
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1644511149
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1644511149
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1644511149
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1644511149
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1644511149
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1644511149
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1644511149
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1644511149
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1644511149
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1644511149
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1644511149
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1644511149
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1644511149
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1644511149
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1644511149
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1644511149
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1644511149
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1644511149
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1644511149
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1644511149
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1644511149
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1644511149
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1644511149
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1644511149
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1644511149
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1644511149
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1644511149
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1644511149
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1644511149
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1644511149
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1644511149
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1644511149
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1644511149
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1644511149
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1644511149
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1644511149
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1644511149
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1644511149
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1644511149
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1644511149
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1644511149
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1644511149
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1644511149
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1644511149
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1644511149
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1644511149
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1644511149
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1644511149
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1644511149
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1644511149
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1644511149
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1644511149
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1644511149
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1644511149
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1644511149
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1644511149
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1644511149
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1644511149
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1644511149
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1644511149
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1644511149
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1644511149
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1644511149
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1644511149
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1644511149
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1644511149
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1644511149
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1644511149
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1644511149
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1644511149
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1644511149
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1644511149
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1644511149
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1644511149
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1644511149
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1644511149
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1644511149
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1644511149
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1644511149
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1644511149
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1644511149
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1644511149
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1644511149
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1644511149
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1644511149
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1644511149
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1644511149
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1644511149
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1644511149
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1644511149
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1644511149
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1644511149
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1644511149
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1644511149
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1644511149
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1644511149
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1644511149
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1644511149
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1644511149
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1644511149
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1644511149
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1644511149
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1644511149
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1644511149
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1644511149
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1644511149
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1644511149
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1644511149
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1644511149
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1644511149
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1644511149
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1644511149
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1644511149
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1644511149
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1644511149
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1644511149
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1644511149
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1644511149
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1644511149
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1644511149
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1644511149
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1644511149
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1644511149
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1644511149
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1644511149
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1644511149
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1644511149
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1644511149
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1644511149
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1644511149
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1644511149
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1644511149
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1644511149
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1644511149
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1644511149
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1644511149
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1644511149
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1644511149
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1644511149
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1644511149
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1644511149
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1644511149
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1644511149
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1644511149
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1644511149
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1644511149
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1644511149
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1644511149
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1644511149
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1644511149
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1644511149
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1644511149
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1644511149
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1644511149
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1644511149
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1644511149
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1644511149
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1644511149
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1644511149
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1644511149
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1644511149
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1644511149
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1644511149
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1644511149
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1644511149
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1644511149
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1644511149
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1644511149
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1644511149
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1644511149
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1644511149
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1644511149
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1644511149
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1644511149
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1644511149
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1644511149
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1644511149
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1644511149
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1644511149
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1644511149
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1644511149
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1644511149
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1644511149
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1644511149
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1644511149
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1644511149
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1644511149
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1644511149
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1644511149
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1644511149
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1644511149
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1644511149
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1644511149
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1644511149
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1644511149
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1644511149
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1644511149
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1644511149
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1644511149
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1644511149
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1644511149
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1644511149
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1644511149
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1644511149
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1644511149
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1644511149
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1644511149
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1644511149
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1644511149
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1644511149
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1644511149
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1644511149
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1644511149
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1644511149
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1644511149
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1644511149
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1644511149
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1644511149
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1644511149
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1644511149
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1644511149
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1644511149
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1644511149
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1644511149
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1644511149
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1644511149
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1644511149
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1644511149
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1644511149
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1644511149
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1644511149
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1644511149
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1644511149
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1644511149
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1644511149
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1644511149
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1644511149
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1644511149
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1644511149
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1644511149
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1644511149
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1644511149
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1644511149
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1644511149
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1644511149
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1644511149
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1644511149
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1644511149
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1644511149
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1644511149
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1644511149
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1644511149
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1644511149
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1644511149
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1644511149
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1644511149
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1644511149
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1644511149
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1644511149
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1644511149
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1644511149
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1644511149
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1644511149
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1644511149
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1644511149
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1644511149
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1644511149
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1644511149
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1644511149
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1644511149
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1644511149
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1644511149
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1644511149
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1644511149
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1644511149
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1644511149
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1644511149
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1644511149
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1644511149
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1644511149
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1644511149
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1644511149
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1644511149
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1644511149
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1644511149
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1644511149
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1644511149
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1644511149
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1644511149
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1644511149
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1644511149
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1644511149
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1644511149
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1644511149
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1644511149
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1644511149
transform 1 0 60352 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1644511149
transform 1 0 65504 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1644511149
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1644511149
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1644511149
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1644511149
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1644511149
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1644511149
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1644511149
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1644511149
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1644511149
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1644511149
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1644511149
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1644511149
transform 1 0 62928 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1644511149
transform 1 0 68080 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1644511149
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1644511149
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1644511149
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1644511149
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1644511149
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1644511149
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1644511149
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1644511149
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1644511149
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1644511149
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1644511149
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1644511149
transform 1 0 60352 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1644511149
transform 1 0 65504 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1644511149
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1644511149
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1644511149
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1644511149
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1644511149
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1644511149
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1644511149
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1644511149
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1644511149
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1644511149
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1644511149
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1644511149
transform 1 0 62928 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1644511149
transform 1 0 68080 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1644511149
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1644511149
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1644511149
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1644511149
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1644511149
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1644511149
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1644511149
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1644511149
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1644511149
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1644511149
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1644511149
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1644511149
transform 1 0 60352 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1644511149
transform 1 0 65504 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1644511149
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1644511149
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1644511149
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1644511149
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1644511149
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1644511149
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1644511149
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1644511149
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1660
timestamp 1644511149
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1661
timestamp 1644511149
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1662
timestamp 1644511149
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1663
timestamp 1644511149
transform 1 0 62928 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1664
timestamp 1644511149
transform 1 0 68080 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1665
timestamp 1644511149
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1666
timestamp 1644511149
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1667
timestamp 1644511149
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1668
timestamp 1644511149
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1669
timestamp 1644511149
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1670
timestamp 1644511149
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1671
timestamp 1644511149
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1672
timestamp 1644511149
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1673
timestamp 1644511149
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1674
timestamp 1644511149
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1675
timestamp 1644511149
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1676
timestamp 1644511149
transform 1 0 60352 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1677
timestamp 1644511149
transform 1 0 65504 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1678
timestamp 1644511149
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1679
timestamp 1644511149
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1680
timestamp 1644511149
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1681
timestamp 1644511149
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1682
timestamp 1644511149
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1683
timestamp 1644511149
transform 1 0 32016 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1684
timestamp 1644511149
transform 1 0 37168 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1685
timestamp 1644511149
transform 1 0 42320 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1686
timestamp 1644511149
transform 1 0 47472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1687
timestamp 1644511149
transform 1 0 52624 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1688
timestamp 1644511149
transform 1 0 57776 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1689
timestamp 1644511149
transform 1 0 62928 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1690
timestamp 1644511149
transform 1 0 68080 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1691
timestamp 1644511149
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1692
timestamp 1644511149
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1693
timestamp 1644511149
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1694
timestamp 1644511149
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1695
timestamp 1644511149
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1696
timestamp 1644511149
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1697
timestamp 1644511149
transform 1 0 34592 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1698
timestamp 1644511149
transform 1 0 39744 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1699
timestamp 1644511149
transform 1 0 44896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1700
timestamp 1644511149
transform 1 0 50048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1701
timestamp 1644511149
transform 1 0 55200 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1702
timestamp 1644511149
transform 1 0 60352 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1703
timestamp 1644511149
transform 1 0 65504 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1704
timestamp 1644511149
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1705
timestamp 1644511149
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1706
timestamp 1644511149
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1707
timestamp 1644511149
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1708
timestamp 1644511149
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1709
timestamp 1644511149
transform 1 0 32016 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1710
timestamp 1644511149
transform 1 0 37168 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1711
timestamp 1644511149
transform 1 0 42320 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1712
timestamp 1644511149
transform 1 0 47472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1713
timestamp 1644511149
transform 1 0 52624 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1714
timestamp 1644511149
transform 1 0 57776 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1715
timestamp 1644511149
transform 1 0 62928 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1716
timestamp 1644511149
transform 1 0 68080 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1717
timestamp 1644511149
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1718
timestamp 1644511149
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1719
timestamp 1644511149
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1720
timestamp 1644511149
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1721
timestamp 1644511149
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1722
timestamp 1644511149
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1723
timestamp 1644511149
transform 1 0 34592 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1724
timestamp 1644511149
transform 1 0 39744 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1725
timestamp 1644511149
transform 1 0 44896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1726
timestamp 1644511149
transform 1 0 50048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1727
timestamp 1644511149
transform 1 0 55200 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1728
timestamp 1644511149
transform 1 0 60352 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1729
timestamp 1644511149
transform 1 0 65504 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1730
timestamp 1644511149
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1731
timestamp 1644511149
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1732
timestamp 1644511149
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1733
timestamp 1644511149
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1734
timestamp 1644511149
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1735
timestamp 1644511149
transform 1 0 32016 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1736
timestamp 1644511149
transform 1 0 37168 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1737
timestamp 1644511149
transform 1 0 42320 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1738
timestamp 1644511149
transform 1 0 47472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1739
timestamp 1644511149
transform 1 0 52624 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1740
timestamp 1644511149
transform 1 0 57776 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1741
timestamp 1644511149
transform 1 0 62928 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1742
timestamp 1644511149
transform 1 0 68080 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1743
timestamp 1644511149
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1744
timestamp 1644511149
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1745
timestamp 1644511149
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1746
timestamp 1644511149
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1747
timestamp 1644511149
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1748
timestamp 1644511149
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1749
timestamp 1644511149
transform 1 0 34592 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1750
timestamp 1644511149
transform 1 0 39744 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1751
timestamp 1644511149
transform 1 0 44896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1752
timestamp 1644511149
transform 1 0 50048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1753
timestamp 1644511149
transform 1 0 55200 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1754
timestamp 1644511149
transform 1 0 60352 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1755
timestamp 1644511149
transform 1 0 65504 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1756
timestamp 1644511149
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1757
timestamp 1644511149
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1758
timestamp 1644511149
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1759
timestamp 1644511149
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1760
timestamp 1644511149
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1761
timestamp 1644511149
transform 1 0 32016 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1762
timestamp 1644511149
transform 1 0 37168 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1763
timestamp 1644511149
transform 1 0 42320 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1764
timestamp 1644511149
transform 1 0 47472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1765
timestamp 1644511149
transform 1 0 52624 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1766
timestamp 1644511149
transform 1 0 57776 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1767
timestamp 1644511149
transform 1 0 62928 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1768
timestamp 1644511149
transform 1 0 68080 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1769
timestamp 1644511149
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1770
timestamp 1644511149
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1771
timestamp 1644511149
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1772
timestamp 1644511149
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1773
timestamp 1644511149
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1774
timestamp 1644511149
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1775
timestamp 1644511149
transform 1 0 34592 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1776
timestamp 1644511149
transform 1 0 39744 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1777
timestamp 1644511149
transform 1 0 44896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1778
timestamp 1644511149
transform 1 0 50048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1779
timestamp 1644511149
transform 1 0 55200 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1780
timestamp 1644511149
transform 1 0 60352 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1781
timestamp 1644511149
transform 1 0 65504 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1782
timestamp 1644511149
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1783
timestamp 1644511149
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1784
timestamp 1644511149
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1785
timestamp 1644511149
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1786
timestamp 1644511149
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1787
timestamp 1644511149
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1788
timestamp 1644511149
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1789
timestamp 1644511149
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1790
timestamp 1644511149
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1791
timestamp 1644511149
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1792
timestamp 1644511149
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1793
timestamp 1644511149
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1794
timestamp 1644511149
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1795
timestamp 1644511149
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1796
timestamp 1644511149
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1797
timestamp 1644511149
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1798
timestamp 1644511149
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1799
timestamp 1644511149
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1800
timestamp 1644511149
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1801
timestamp 1644511149
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1802
timestamp 1644511149
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1803
timestamp 1644511149
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1804
timestamp 1644511149
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1805
timestamp 1644511149
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1806
timestamp 1644511149
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1807
timestamp 1644511149
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1808
timestamp 1644511149
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1809
timestamp 1644511149
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1810
timestamp 1644511149
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1811
timestamp 1644511149
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1812
timestamp 1644511149
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1813
timestamp 1644511149
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1814
timestamp 1644511149
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1815
timestamp 1644511149
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1816
timestamp 1644511149
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1817
timestamp 1644511149
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1818
timestamp 1644511149
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1819
timestamp 1644511149
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1820
timestamp 1644511149
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1821
timestamp 1644511149
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1822
timestamp 1644511149
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1823
timestamp 1644511149
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1824
timestamp 1644511149
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1825
timestamp 1644511149
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1826
timestamp 1644511149
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1827
timestamp 1644511149
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1828
timestamp 1644511149
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1829
timestamp 1644511149
transform 1 0 44896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1830
timestamp 1644511149
transform 1 0 50048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1831
timestamp 1644511149
transform 1 0 55200 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1832
timestamp 1644511149
transform 1 0 60352 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1833
timestamp 1644511149
transform 1 0 65504 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1834
timestamp 1644511149
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1835
timestamp 1644511149
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1836
timestamp 1644511149
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1837
timestamp 1644511149
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1838
timestamp 1644511149
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1839
timestamp 1644511149
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1840
timestamp 1644511149
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1841
timestamp 1644511149
transform 1 0 42320 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1842
timestamp 1644511149
transform 1 0 47472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1843
timestamp 1644511149
transform 1 0 52624 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1844
timestamp 1644511149
transform 1 0 57776 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1845
timestamp 1644511149
transform 1 0 62928 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1846
timestamp 1644511149
transform 1 0 68080 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1847
timestamp 1644511149
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1848
timestamp 1644511149
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1849
timestamp 1644511149
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1850
timestamp 1644511149
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1851
timestamp 1644511149
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1852
timestamp 1644511149
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1853
timestamp 1644511149
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1854
timestamp 1644511149
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1855
timestamp 1644511149
transform 1 0 44896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1856
timestamp 1644511149
transform 1 0 50048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1857
timestamp 1644511149
transform 1 0 55200 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1858
timestamp 1644511149
transform 1 0 60352 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1859
timestamp 1644511149
transform 1 0 65504 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1860
timestamp 1644511149
transform 1 0 3680 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1861
timestamp 1644511149
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1862
timestamp 1644511149
transform 1 0 8832 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1863
timestamp 1644511149
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1864
timestamp 1644511149
transform 1 0 13984 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1865
timestamp 1644511149
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1866
timestamp 1644511149
transform 1 0 19136 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1867
timestamp 1644511149
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1868
timestamp 1644511149
transform 1 0 24288 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1869
timestamp 1644511149
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1870
timestamp 1644511149
transform 1 0 29440 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1871
timestamp 1644511149
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1872
timestamp 1644511149
transform 1 0 34592 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1873
timestamp 1644511149
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1874
timestamp 1644511149
transform 1 0 39744 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1875
timestamp 1644511149
transform 1 0 42320 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1876
timestamp 1644511149
transform 1 0 44896 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1877
timestamp 1644511149
transform 1 0 47472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1878
timestamp 1644511149
transform 1 0 50048 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1879
timestamp 1644511149
transform 1 0 52624 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1880
timestamp 1644511149
transform 1 0 55200 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1881
timestamp 1644511149
transform 1 0 57776 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1882
timestamp 1644511149
transform 1 0 60352 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1883
timestamp 1644511149
transform 1 0 62928 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1884
timestamp 1644511149
transform 1 0 65504 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1885
timestamp 1644511149
transform 1 0 68080 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _242_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _243_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33488 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _244_
timestamp 1644511149
transform 1 0 27140 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _245_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1644511149
transform -1 0 12236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1644511149
transform 1 0 28336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1644511149
transform -1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _250_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1644511149
transform 1 0 27876 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1644511149
transform 1 0 59708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1644511149
transform -1 0 23920 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1644511149
transform 1 0 60536 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1644511149
transform 1 0 60444 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _256_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36524 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _257_
timestamp 1644511149
transform -1 0 35972 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1644511149
transform 1 0 50876 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1644511149
transform -1 0 32292 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1644511149
transform 1 0 54096 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1644511149
transform -1 0 32384 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1644511149
transform 1 0 36524 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _263_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36156 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1644511149
transform -1 0 28704 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1644511149
transform -1 0 61364 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1644511149
transform 1 0 61640 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1644511149
transform -1 0 25024 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1644511149
transform 1 0 60996 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _269_
timestamp 1644511149
transform -1 0 35880 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1644511149
transform 1 0 53452 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1644511149
transform 1 0 41308 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1644511149
transform -1 0 24840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1644511149
transform 1 0 50416 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _275_
timestamp 1644511149
transform -1 0 36156 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1644511149
transform 1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1644511149
transform 1 0 47104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1644511149
transform -1 0 10580 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1644511149
transform 1 0 43332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _281_
timestamp 1644511149
transform -1 0 36156 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1644511149
transform 1 0 51428 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1644511149
transform 1 0 54188 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1644511149
transform 1 0 45908 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1644511149
transform -1 0 23736 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1644511149
transform 1 0 26220 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _287_
timestamp 1644511149
transform 1 0 35328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _288_
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1644511149
transform 1 0 51520 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1644511149
transform 1 0 31740 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1644511149
transform 1 0 48576 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1644511149
transform -1 0 26220 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1644511149
transform -1 0 28520 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _294_
timestamp 1644511149
transform -1 0 37168 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1644511149
transform -1 0 9844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1644511149
transform 1 0 44528 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1644511149
transform -1 0 10304 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1644511149
transform -1 0 9752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1644511149
transform 1 0 41492 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _300_
timestamp 1644511149
transform 1 0 38456 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1644511149
transform 1 0 64860 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1644511149
transform -1 0 34960 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1644511149
transform 1 0 64676 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1644511149
transform -1 0 64400 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1644511149
transform 1 0 64768 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _306_
timestamp 1644511149
transform 1 0 37444 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1644511149
transform -1 0 25392 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1644511149
transform 1 0 50692 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1644511149
transform -1 0 22080 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1644511149
transform 1 0 43884 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1644511149
transform 1 0 49036 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _312_
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1644511149
transform 1 0 38180 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1644511149
transform 1 0 44896 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1644511149
transform -1 0 24932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1644511149
transform 1 0 46828 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1644511149
transform -1 0 28060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _318_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33028 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _319_
timestamp 1644511149
transform -1 0 33764 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1644511149
transform 1 0 43976 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1644511149
transform 1 0 8372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1644511149
transform -1 0 9200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1644511149
transform -1 0 8464 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1644511149
transform 1 0 40020 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _325_
timestamp 1644511149
transform 1 0 39652 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1644511149
transform 1 0 63940 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1644511149
transform -1 0 63756 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1644511149
transform -1 0 37536 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1644511149
transform 1 0 64584 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1644511149
transform -1 0 56304 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _331_
timestamp 1644511149
transform 1 0 38180 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1644511149
transform 1 0 56764 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1644511149
transform 1 0 35696 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1644511149
transform 1 0 58788 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1644511149
transform -1 0 34776 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1644511149
transform 1 0 58144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _337_
timestamp 1644511149
transform -1 0 33580 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1644511149
transform 1 0 16836 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1644511149
transform -1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1644511149
transform 1 0 14996 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1644511149
transform -1 0 13156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _343_
timestamp 1644511149
transform -1 0 39284 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1644511149
transform 1 0 61640 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1644511149
transform 1 0 62192 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1644511149
transform -1 0 30820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1644511149
transform -1 0 28244 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1644511149
transform 1 0 62008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _349_
timestamp 1644511149
transform 1 0 32292 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1644511149
transform -1 0 20148 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1644511149
transform 1 0 43332 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1644511149
transform -1 0 20332 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1644511149
transform -1 0 19688 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _355_
timestamp 1644511149
transform 1 0 33948 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1644511149
transform -1 0 34960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1644511149
transform -1 0 34960 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1644511149
transform 1 0 35604 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1644511149
transform 1 0 51612 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1644511149
transform 1 0 49128 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _361_
timestamp 1644511149
transform 1 0 33856 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1644511149
transform 1 0 40756 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1644511149
transform 1 0 56212 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1644511149
transform 1 0 57224 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1644511149
transform -1 0 33764 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1644511149
transform -1 0 56580 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _367_
timestamp 1644511149
transform -1 0 33028 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1644511149
transform -1 0 6624 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1644511149
transform 1 0 35144 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1644511149
transform -1 0 14352 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1644511149
transform -1 0 6624 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1644511149
transform -1 0 6624 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1644511149
transform -1 0 27232 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1644511149
transform 1 0 36156 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _376__2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _377__3
timestamp 1644511149
transform -1 0 12052 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _378__4
timestamp 1644511149
transform -1 0 29808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _379__5
timestamp 1644511149
transform 1 0 10488 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _380__6
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _381__7
timestamp 1644511149
transform 1 0 28520 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _382__8
timestamp 1644511149
transform 1 0 59984 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _383__9
timestamp 1644511149
transform 1 0 23000 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _384__10
timestamp 1644511149
transform -1 0 61272 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _385__11
timestamp 1644511149
transform -1 0 60720 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _386__12
timestamp 1644511149
transform -1 0 51428 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _387__13
timestamp 1644511149
transform -1 0 32936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _388__14
timestamp 1644511149
transform 1 0 54556 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _389__15
timestamp 1644511149
transform 1 0 31004 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _390__16
timestamp 1644511149
transform 1 0 36892 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _391__17
timestamp 1644511149
transform -1 0 28428 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _392__18
timestamp 1644511149
transform -1 0 61456 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _393__19
timestamp 1644511149
transform -1 0 62192 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _394__20
timestamp 1644511149
transform 1 0 24288 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _395__21
timestamp 1644511149
transform -1 0 61916 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _396__22
timestamp 1644511149
transform -1 0 26496 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _397__23
timestamp 1644511149
transform -1 0 54464 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _398__24
timestamp 1644511149
transform -1 0 42688 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _399__25
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _400__26
timestamp 1644511149
transform 1 0 49680 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _401__27
timestamp 1644511149
transform -1 0 12236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _402__28
timestamp 1644511149
transform -1 0 48116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _403__29
timestamp 1644511149
transform -1 0 10120 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _404__30
timestamp 1644511149
transform -1 0 43792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _405__31
timestamp 1644511149
transform 1 0 10672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _406__32
timestamp 1644511149
transform 1 0 50784 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _407__33
timestamp 1644511149
transform -1 0 55568 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _408__34
timestamp 1644511149
transform -1 0 37628 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _409__35
timestamp 1644511149
transform -1 0 46184 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _410__36
timestamp 1644511149
transform 1 0 22816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _411__37
timestamp 1644511149
transform 1 0 26312 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _412__38
timestamp 1644511149
transform -1 0 52992 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _413__39
timestamp 1644511149
transform 1 0 31372 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _414__40
timestamp 1644511149
transform 1 0 48484 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _415__41
timestamp 1644511149
transform 1 0 25300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _416__42
timestamp 1644511149
transform -1 0 28336 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _417__43
timestamp 1644511149
transform -1 0 9568 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _418__44
timestamp 1644511149
transform -1 0 45632 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _419__45
timestamp 1644511149
transform 1 0 9384 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _420__46
timestamp 1644511149
transform -1 0 9292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _421__47
timestamp 1644511149
transform -1 0 42688 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _422__48
timestamp 1644511149
transform -1 0 65872 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _423__49
timestamp 1644511149
transform 1 0 33580 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _424__50
timestamp 1644511149
transform -1 0 65872 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _425__51
timestamp 1644511149
transform -1 0 64308 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _426__52
timestamp 1644511149
transform 1 0 65412 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _427__53
timestamp 1644511149
transform -1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _428__54
timestamp 1644511149
transform -1 0 51336 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _429__55
timestamp 1644511149
transform 1 0 20792 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _430__56
timestamp 1644511149
transform -1 0 45264 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _431__57
timestamp 1644511149
transform -1 0 49496 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _432__58
timestamp 1644511149
transform -1 0 39100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _433__59
timestamp 1644511149
transform -1 0 45356 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _434__60
timestamp 1644511149
transform 1 0 24196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _435__61
timestamp 1644511149
transform 1 0 46828 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _436__62
timestamp 1644511149
transform -1 0 27784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _437__63
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _438__64
timestamp 1644511149
transform 1 0 8096 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _439__65
timestamp 1644511149
transform -1 0 9200 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _440__66
timestamp 1644511149
transform -1 0 8096 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _441__67
timestamp 1644511149
transform -1 0 40480 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _442__68
timestamp 1644511149
transform 1 0 63296 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _443__69
timestamp 1644511149
transform -1 0 63940 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _444__70
timestamp 1644511149
transform 1 0 36340 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _445__71
timestamp 1644511149
transform -1 0 65872 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _446__72
timestamp 1644511149
transform -1 0 37536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _447__73
timestamp 1644511149
transform -1 0 56120 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _448__74
timestamp 1644511149
transform -1 0 58144 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _449__75
timestamp 1644511149
transform -1 0 36616 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _450__76
timestamp 1644511149
transform -1 0 59708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _451__77
timestamp 1644511149
transform 1 0 33948 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _452__78
timestamp 1644511149
transform -1 0 58512 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _453__79
timestamp 1644511149
transform -1 0 17112 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _454__80
timestamp 1644511149
transform -1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _455__81
timestamp 1644511149
transform -1 0 15272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _456__82
timestamp 1644511149
transform -1 0 12604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _457__83
timestamp 1644511149
transform -1 0 33304 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _458__84
timestamp 1644511149
transform -1 0 62100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _459__85
timestamp 1644511149
transform 1 0 62468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _460__86
timestamp 1644511149
transform 1 0 31188 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _461__87
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _462__88
timestamp 1644511149
transform 1 0 62652 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _463__89
timestamp 1644511149
transform -1 0 19780 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _464__90
timestamp 1644511149
transform -1 0 44252 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _465__91
timestamp 1644511149
transform -1 0 20056 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _466__92
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _467__93
timestamp 1644511149
transform 1 0 18768 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _468__94
timestamp 1644511149
transform -1 0 34040 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _469__95
timestamp 1644511149
transform -1 0 34960 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _470__96
timestamp 1644511149
transform -1 0 35880 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _471__97
timestamp 1644511149
transform 1 0 51980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _472__98
timestamp 1644511149
transform -1 0 49496 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _473__99
timestamp 1644511149
transform -1 0 41032 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _474__100
timestamp 1644511149
transform -1 0 56672 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _475__101
timestamp 1644511149
transform -1 0 58236 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _476__102
timestamp 1644511149
transform -1 0 33212 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _477__103
timestamp 1644511149
transform -1 0 56672 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _478__104
timestamp 1644511149
transform 1 0 6164 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _479__105
timestamp 1644511149
transform -1 0 36064 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _480__106
timestamp 1644511149
transform 1 0 13248 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _481__107
timestamp 1644511149
transform -1 0 5704 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _482__108
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _483__109
timestamp 1644511149
transform 1 0 25944 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _484_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13616 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _485_
timestamp 1644511149
transform 1 0 11684 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _486_
timestamp 1644511149
transform 1 0 28980 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _487_
timestamp 1644511149
transform -1 0 12328 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _488_
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _489_
timestamp 1644511149
transform -1 0 29072 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _490_
timestamp 1644511149
transform 1 0 60444 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _491_
timestamp 1644511149
transform 1 0 23092 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _492_
timestamp 1644511149
transform 1 0 60628 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _493_
timestamp 1644511149
transform 1 0 60260 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _494_
timestamp 1644511149
transform 1 0 51060 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _495_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _496_
timestamp 1644511149
transform 1 0 55292 0 1 60928
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _497_
timestamp 1644511149
transform -1 0 32844 0 1 62016
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _498_
timestamp 1644511149
transform 1 0 37260 0 -1 62016
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _499_
timestamp 1644511149
transform 1 0 28152 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _500_
timestamp 1644511149
transform 1 0 60628 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _501_
timestamp 1644511149
transform 1 0 61916 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _502_
timestamp 1644511149
transform 1 0 24380 0 1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _503_
timestamp 1644511149
transform 1 0 61640 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _504_
timestamp 1644511149
transform 1 0 26128 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _505_
timestamp 1644511149
transform 1 0 54096 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _506_
timestamp 1644511149
transform 1 0 41952 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _507_
timestamp 1644511149
transform 1 0 24104 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _508_
timestamp 1644511149
transform 1 0 50324 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _509_
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _510_
timestamp 1644511149
transform 1 0 47748 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _511_
timestamp 1644511149
transform 1 0 9752 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _512_
timestamp 1644511149
transform 1 0 43424 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _513_
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _514_
timestamp 1644511149
transform 1 0 51520 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _515_
timestamp 1644511149
transform 1 0 54832 0 -1 59840
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _516_
timestamp 1644511149
transform 1 0 37352 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _517_
timestamp 1644511149
transform 1 0 45816 0 1 60928
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _518_
timestamp 1644511149
transform 1 0 23000 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _519_
timestamp 1644511149
transform 1 0 26956 0 -1 59840
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _520_
timestamp 1644511149
transform 1 0 52164 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _521_
timestamp 1644511149
transform 1 0 32108 0 -1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _522_
timestamp 1644511149
transform 1 0 48668 0 -1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _523_
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _524_
timestamp 1644511149
transform 1 0 27968 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _525_
timestamp 1644511149
transform 1 0 9292 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _526_
timestamp 1644511149
transform 1 0 45172 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _527_
timestamp 1644511149
transform 1 0 9752 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _528_
timestamp 1644511149
transform 1 0 9016 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _529_
timestamp 1644511149
transform 1 0 41676 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _530_
timestamp 1644511149
transform 1 0 64952 0 -1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _531_
timestamp 1644511149
transform -1 0 35420 0 -1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _532_
timestamp 1644511149
transform 1 0 65320 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _533_
timestamp 1644511149
transform 1 0 63940 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _534_
timestamp 1644511149
transform 1 0 65596 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _535_
timestamp 1644511149
transform 1 0 24840 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _536_
timestamp 1644511149
transform 1 0 50968 0 1 51136
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _537_
timestamp 1644511149
transform -1 0 22724 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _538_
timestamp 1644511149
transform 1 0 44528 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _539_
timestamp 1644511149
transform 1 0 49128 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _540_
timestamp 1644511149
transform 1 0 38088 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _541_
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _542_
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _543_
timestamp 1644511149
transform 1 0 47564 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _544_
timestamp 1644511149
transform 1 0 27508 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _545_
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _546_
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _547_
timestamp 1644511149
transform 1 0 8648 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _548_
timestamp 1644511149
transform 1 0 7728 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _549_
timestamp 1644511149
transform 1 0 40020 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _550_
timestamp 1644511149
transform 1 0 64032 0 -1 57664
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _551_
timestamp 1644511149
transform 1 0 63204 0 1 54400
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _552_
timestamp 1644511149
transform -1 0 38180 0 1 57664
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _553_
timestamp 1644511149
transform 1 0 64308 0 -1 58752
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _554_
timestamp 1644511149
transform 1 0 36800 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _555_
timestamp 1644511149
transform 1 0 55476 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _556_
timestamp 1644511149
transform 1 0 57408 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _557_
timestamp 1644511149
transform 1 0 35604 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _558_
timestamp 1644511149
transform 1 0 59156 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _559_
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _560_
timestamp 1644511149
transform 1 0 58052 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _561_
timestamp 1644511149
transform 1 0 16744 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _562_
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _563_
timestamp 1644511149
transform 1 0 14904 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _564_
timestamp 1644511149
transform 1 0 12328 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _565_
timestamp 1644511149
transform 1 0 32936 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _566_
timestamp 1644511149
transform 1 0 61732 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _567_
timestamp 1644511149
transform 1 0 63020 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _568_
timestamp 1644511149
transform -1 0 32200 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _569_
timestamp 1644511149
transform 1 0 27508 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _570_
timestamp 1644511149
transform 1 0 63020 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _571_
timestamp 1644511149
transform 1 0 19412 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _572_
timestamp 1644511149
transform 1 0 43608 0 -1 63104
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _573_
timestamp 1644511149
transform 1 0 19412 0 -1 64192
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _574_
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _575_
timestamp 1644511149
transform 1 0 19320 0 1 63104
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _576_
timestamp 1644511149
transform 1 0 33764 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _577_
timestamp 1644511149
transform 1 0 34224 0 -1 57664
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _578_
timestamp 1644511149
transform 1 0 35512 0 1 58752
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _579_
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _580_
timestamp 1644511149
transform 1 0 49220 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _581_
timestamp 1644511149
transform 1 0 40664 0 1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _582_
timestamp 1644511149
transform 1 0 56304 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _583_
timestamp 1644511149
transform 1 0 57868 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _584_
timestamp 1644511149
transform 1 0 32936 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _585_
timestamp 1644511149
transform 1 0 55752 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _586_
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _587_
timestamp 1644511149
transform 1 0 35512 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _588_
timestamp 1644511149
transform 1 0 13892 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _589_
timestamp 1644511149
transform 1 0 5428 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _590_
timestamp 1644511149
transform -1 0 7636 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _591_
timestamp 1644511149
transform -1 0 27784 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1644511149
transform 1 0 1380 0 -1 66368
box -38 -48 590 592
<< labels >>
rlabel metal3 s 0 65908 800 66148 6 active
port 0 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 38630 71200 38742 72000 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 71348 800 71588 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 69200 60468 70000 60708 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 25750 71200 25862 72000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 69200 63188 70000 63428 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 69200 6748 70000 6988 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 13514 71200 13626 72000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 16090 71200 16202 72000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 61170 0 61282 800 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 69200 23748 70000 23988 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 12226 71200 12338 72000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 8362 71200 8474 72000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 53442 0 53554 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 52154 0 52266 800 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 69200 16268 70000 16508 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 69542 71200 69654 72000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 69200 29188 70000 29428 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 63188 800 63428 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 52798 71200 52910 72000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 60526 71200 60638 72000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 69200 45508 70000 45748 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 61814 71200 61926 72000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 39918 71200 40030 72000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 69200 44148 70000 44388 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 69200 68628 70000 68868 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 0 43468 800 43708 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 69200 48228 70000 48468 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 10938 71200 11050 72000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 io_oeb[0]
port 39 nsew signal bidirectional
rlabel metal3 s 0 24428 800 24668 6 io_oeb[10]
port 40 nsew signal bidirectional
rlabel metal3 s 69200 41428 70000 41668 6 io_oeb[11]
port 41 nsew signal bidirectional
rlabel metal3 s 69200 21708 70000 21948 6 io_oeb[12]
port 42 nsew signal bidirectional
rlabel metal3 s 69200 20348 70000 20588 6 io_oeb[13]
port 43 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 io_oeb[14]
port 44 nsew signal bidirectional
rlabel metal2 s 18666 71200 18778 72000 6 io_oeb[15]
port 45 nsew signal bidirectional
rlabel metal3 s 69200 4028 70000 4268 6 io_oeb[16]
port 46 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 io_oeb[17]
port 47 nsew signal bidirectional
rlabel metal2 s 50222 71200 50334 72000 6 io_oeb[18]
port 48 nsew signal bidirectional
rlabel metal2 s 19954 71200 20066 72000 6 io_oeb[19]
port 49 nsew signal bidirectional
rlabel metal2 s 56018 0 56130 800 6 io_oeb[1]
port 50 nsew signal bidirectional
rlabel metal3 s 69200 31908 70000 32148 6 io_oeb[20]
port 51 nsew signal bidirectional
rlabel metal2 s 1922 71200 2034 72000 6 io_oeb[21]
port 52 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 io_oeb[22]
port 53 nsew signal bidirectional
rlabel metal2 s 34766 71200 34878 72000 6 io_oeb[23]
port 54 nsew signal bidirectional
rlabel metal2 s 36054 71200 36166 72000 6 io_oeb[24]
port 55 nsew signal bidirectional
rlabel metal2 s 67610 0 67722 800 6 io_oeb[25]
port 56 nsew signal bidirectional
rlabel metal3 s 69200 56388 70000 56628 6 io_oeb[26]
port 57 nsew signal bidirectional
rlabel metal2 s 41206 71200 41318 72000 6 io_oeb[27]
port 58 nsew signal bidirectional
rlabel metal2 s 59882 0 59994 800 6 io_oeb[28]
port 59 nsew signal bidirectional
rlabel metal3 s 69200 46868 70000 47108 6 io_oeb[29]
port 60 nsew signal bidirectional
rlabel metal2 s 57950 71200 58062 72000 6 io_oeb[2]
port 61 nsew signal bidirectional
rlabel metal2 s 3210 71200 3322 72000 6 io_oeb[30]
port 62 nsew signal bidirectional
rlabel metal2 s 58594 0 58706 800 6 io_oeb[31]
port 63 nsew signal bidirectional
rlabel metal3 s 0 35308 800 35548 6 io_oeb[32]
port 64 nsew signal bidirectional
rlabel metal2 s 68898 0 69010 800 6 io_oeb[33]
port 65 nsew signal bidirectional
rlabel metal2 s 14802 71200 14914 72000 6 io_oeb[34]
port 66 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 io_oeb[35]
port 67 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 io_oeb[36]
port 68 nsew signal bidirectional
rlabel metal3 s 0 25788 800 26028 6 io_oeb[37]
port 69 nsew signal bidirectional
rlabel metal2 s 36054 0 36166 800 6 io_oeb[3]
port 70 nsew signal bidirectional
rlabel metal3 s 69200 1308 70000 1548 6 io_oeb[4]
port 71 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 io_oeb[5]
port 72 nsew signal bidirectional
rlabel metal3 s 69200 26468 70000 26708 6 io_oeb[6]
port 73 nsew signal bidirectional
rlabel metal2 s 17378 71200 17490 72000 6 io_oeb[7]
port 74 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 io_oeb[8]
port 75 nsew signal bidirectional
rlabel metal2 s 15446 0 15558 800 6 io_oeb[9]
port 76 nsew signal bidirectional
rlabel metal3 s 69200 67268 70000 67508 6 io_out[0]
port 77 nsew signal bidirectional
rlabel metal3 s 69200 40068 70000 40308 6 io_out[10]
port 78 nsew signal bidirectional
rlabel metal3 s 0 4028 800 4268 6 io_out[11]
port 79 nsew signal bidirectional
rlabel metal3 s 0 10828 800 11068 6 io_out[12]
port 80 nsew signal bidirectional
rlabel metal2 s 57306 0 57418 800 6 io_out[13]
port 81 nsew signal bidirectional
rlabel metal3 s 69200 57748 70000 57988 6 io_out[14]
port 82 nsew signal bidirectional
rlabel metal3 s 0 59108 800 59348 6 io_out[15]
port 83 nsew signal bidirectional
rlabel metal3 s 69200 38708 70000 38948 6 io_out[16]
port 84 nsew signal bidirectional
rlabel metal2 s 64390 71200 64502 72000 6 io_out[17]
port 85 nsew signal bidirectional
rlabel metal2 s 66322 0 66434 800 6 io_out[18]
port 86 nsew signal bidirectional
rlabel metal3 s 0 33948 800 34188 6 io_out[19]
port 87 nsew signal bidirectional
rlabel metal2 s 46358 71200 46470 72000 6 io_out[1]
port 88 nsew signal bidirectional
rlabel metal2 s 56662 71200 56774 72000 6 io_out[20]
port 89 nsew signal bidirectional
rlabel metal3 s 0 57748 800 57988 6 io_out[21]
port 90 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 io_out[22]
port 91 nsew signal bidirectional
rlabel metal3 s 69200 33268 70000 33508 6 io_out[23]
port 92 nsew signal bidirectional
rlabel metal2 s 38630 0 38742 800 6 io_out[24]
port 93 nsew signal bidirectional
rlabel metal2 s 51510 71200 51622 72000 6 io_out[25]
port 94 nsew signal bidirectional
rlabel metal3 s 0 8108 800 8348 6 io_out[26]
port 95 nsew signal bidirectional
rlabel metal2 s 54086 71200 54198 72000 6 io_out[27]
port 96 nsew signal bidirectional
rlabel metal2 s 24462 0 24574 800 6 io_out[28]
port 97 nsew signal bidirectional
rlabel metal3 s 69200 2668 70000 2908 6 io_out[29]
port 98 nsew signal bidirectional
rlabel metal2 s 10294 0 10406 800 6 io_out[2]
port 99 nsew signal bidirectional
rlabel metal3 s 0 9468 800 9708 6 io_out[30]
port 100 nsew signal bidirectional
rlabel metal3 s 0 20348 800 20588 6 io_out[31]
port 101 nsew signal bidirectional
rlabel metal3 s 0 67268 800 67508 6 io_out[32]
port 102 nsew signal bidirectional
rlabel metal3 s 69200 10828 70000 11068 6 io_out[33]
port 103 nsew signal bidirectional
rlabel metal3 s 69200 59108 70000 59348 6 io_out[34]
port 104 nsew signal bidirectional
rlabel metal3 s 69200 55028 70000 55268 6 io_out[35]
port 105 nsew signal bidirectional
rlabel metal2 s 21242 71200 21354 72000 6 io_out[36]
port 106 nsew signal bidirectional
rlabel metal3 s 69200 64548 70000 64788 6 io_out[37]
port 107 nsew signal bidirectional
rlabel metal3 s 0 61828 800 62068 6 io_out[3]
port 108 nsew signal bidirectional
rlabel metal3 s 69200 42788 70000 43028 6 io_out[4]
port 109 nsew signal bidirectional
rlabel metal2 s 32190 71200 32302 72000 6 io_out[5]
port 110 nsew signal bidirectional
rlabel metal2 s 66966 71200 67078 72000 6 io_out[6]
port 111 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 io_out[7]
port 112 nsew signal bidirectional
rlabel metal2 s 27038 0 27150 800 6 io_out[8]
port 113 nsew signal bidirectional
rlabel metal3 s 0 21708 800 21948 6 io_out[9]
port 114 nsew signal bidirectional
rlabel metal3 s 69200 12188 70000 12428 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 30902 0 31014 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal3 s 69200 9468 70000 9708 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal3 s 0 53668 800 53908 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 18988 800 19228 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 22530 71200 22642 72000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 43782 71200 43894 72000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 33478 71200 33590 72000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal2 s 62458 0 62570 800 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 24462 71200 24574 72000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal3 s 0 52308 800 52548 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 68254 71200 68366 72000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal3 s 69200 13548 70000 13788 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 1308 800 1548 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal3 s 0 55028 800 55268 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal3 s 69200 5388 70000 5628 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal2 s 634 71200 746 72000 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal2 s 54730 0 54842 800 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 59238 71200 59350 72000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 69200 35988 70000 36228 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 27038 71200 27150 72000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 28326 71200 28438 72000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_data_out[0]
port 147 nsew signal bidirectional
rlabel metal3 s 69200 17628 70000 17868 6 la1_data_out[10]
port 148 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la1_data_out[11]
port 149 nsew signal bidirectional
rlabel metal3 s 69200 65908 70000 66148 6 la1_data_out[12]
port 150 nsew signal bidirectional
rlabel metal2 s 5786 71200 5898 72000 6 la1_data_out[13]
port 151 nsew signal bidirectional
rlabel metal2 s 37342 71200 37454 72000 6 la1_data_out[14]
port 152 nsew signal bidirectional
rlabel metal3 s 0 2668 800 2908 6 la1_data_out[15]
port 153 nsew signal bidirectional
rlabel metal3 s 69200 25108 70000 25348 6 la1_data_out[16]
port 154 nsew signal bidirectional
rlabel metal3 s 69200 52308 70000 52548 6 la1_data_out[17]
port 155 nsew signal bidirectional
rlabel metal2 s 7074 71200 7186 72000 6 la1_data_out[18]
port 156 nsew signal bidirectional
rlabel metal3 s 69200 37348 70000 37588 6 la1_data_out[19]
port 157 nsew signal bidirectional
rlabel metal3 s 0 64548 800 64788 6 la1_data_out[1]
port 158 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la1_data_out[20]
port 159 nsew signal bidirectional
rlabel metal3 s 69200 61828 70000 62068 6 la1_data_out[21]
port 160 nsew signal bidirectional
rlabel metal2 s 42494 71200 42606 72000 6 la1_data_out[22]
port 161 nsew signal bidirectional
rlabel metal2 s 18022 0 18134 800 6 la1_data_out[23]
port 162 nsew signal bidirectional
rlabel metal3 s 69200 27828 70000 28068 6 la1_data_out[24]
port 163 nsew signal bidirectional
rlabel metal3 s 0 5388 800 5628 6 la1_data_out[25]
port 164 nsew signal bidirectional
rlabel metal3 s 69200 8108 70000 8348 6 la1_data_out[26]
port 165 nsew signal bidirectional
rlabel metal3 s 0 68628 800 68868 6 la1_data_out[27]
port 166 nsew signal bidirectional
rlabel metal2 s 63746 0 63858 800 6 la1_data_out[28]
port 167 nsew signal bidirectional
rlabel metal2 s 9006 0 9118 800 6 la1_data_out[29]
port 168 nsew signal bidirectional
rlabel metal2 s 29614 0 29726 800 6 la1_data_out[2]
port 169 nsew signal bidirectional
rlabel metal3 s 69200 18988 70000 19228 6 la1_data_out[30]
port 170 nsew signal bidirectional
rlabel metal3 s 69200 69988 70000 70228 6 la1_data_out[31]
port 171 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la1_data_out[3]
port 172 nsew signal bidirectional
rlabel metal2 s 65034 0 65146 800 6 la1_data_out[4]
port 173 nsew signal bidirectional
rlabel metal2 s 5142 0 5254 800 6 la1_data_out[5]
port 174 nsew signal bidirectional
rlabel metal3 s 69200 30548 70000 30788 6 la1_data_out[6]
port 175 nsew signal bidirectional
rlabel metal2 s 1278 0 1390 800 6 la1_data_out[7]
port 176 nsew signal bidirectional
rlabel metal3 s 69200 53668 70000 53908 6 la1_data_out[8]
port 177 nsew signal bidirectional
rlabel metal2 s 65678 71200 65790 72000 6 la1_data_out[9]
port 178 nsew signal bidirectional
rlabel metal3 s 69200 -52 70000 188 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 63102 71200 63214 72000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 42494 0 42606 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 50866 0 50978 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal3 s 0 50948 800 51188 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal2 s 4498 71200 4610 72000 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 30902 71200 31014 72000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 3854 0 3966 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 45070 71200 45182 72000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 29614 71200 29726 72000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 55374 71200 55486 72000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal3 s 69200 14908 70000 15148 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal3 s 0 56388 800 56628 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 69200 50948 70000 51188 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 69200 49588 70000 49828 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 48934 71200 49046 72000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 47646 71200 47758 72000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal3 s 0 69988 800 70228 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal2 s 9650 71200 9762 72000 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal3 s 0 60468 800 60708 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 4208 2128 4528 69680 6 vccd1
port 211 nsew power input
rlabel metal4 s 34928 2128 35248 69680 6 vccd1
port 211 nsew power input
rlabel metal4 s 65648 2128 65968 69680 6 vccd1
port 211 nsew power input
rlabel metal4 s 19568 2128 19888 69680 6 vssd1
port 212 nsew ground input
rlabel metal4 s 50288 2128 50608 69680 6 vssd1
port 212 nsew ground input
rlabel metal3 s 69200 34628 70000 34868 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 72000
<< end >>
