* NGSPICE file created from wrapped_etpu.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

.subckt wrapped_etpu active vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_159__58 vssd1 vssd1 vccd1 vccd1 _159__58/HI _192_/A sky130_fd_sc_hd__conb_1
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_200_ _200_/A _121_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__ebufn_8
XFILLER_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_131_ _131_/A _131_/B _131_/C _131_/D vssd1 vssd1 vccd1 vccd1 _134_/B sky130_fd_sc_hd__or4_1
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_143__42 vssd1 vssd1 vccd1 vccd1 _143__42/HI _176_/A sky130_fd_sc_hd__conb_1
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_114_ _115_/A vssd1 vssd1 vccd1 vccd1 _114_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_5 _131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_130_ _130_/A _130_/B _130_/C _130_/D vssd1 vssd1 vccd1 vccd1 _134_/A sky130_fd_sc_hd__or4_1
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_113_ _115_/A vssd1 vssd1 vccd1 vccd1 _113_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_6 _131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_164__63 vssd1 vssd1 vccd1 vccd1 _164__63/HI _197_/A sky130_fd_sc_hd__conb_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_189_ _189_/A _108_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__ebufn_8
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_112_ _115_/A vssd1 vssd1 vccd1 vccd1 _112_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_7 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_188_ _188_/A _107_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__ebufn_8
XFILLER_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_111_ _115_/A vssd1 vssd1 vccd1 vccd1 _111_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_8 _130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_155__54 vssd1 vssd1 vccd1 vccd1 _155__54/HI _188_/A sky130_fd_sc_hd__conb_1
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_187_ _187_/A _106_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__ebufn_8
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_110_ _116_/A vssd1 vssd1 vccd1 vccd1 _115_/A sky130_fd_sc_hd__buf_6
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_9 _132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_186_ _186_/A _105_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__ebufn_8
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_140__39 vssd1 vssd1 vccd1 vccd1 _140__39/HI _173_/A sky130_fd_sc_hd__conb_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_169_ _169_/A _129_/A vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__ebufn_8
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_146__45 vssd1 vssd1 vccd1 vccd1 _146__45/HI _179_/A sky130_fd_sc_hd__conb_1
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_185_ _185_/A _103_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__ebufn_8
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_099_ _103_/A vssd1 vssd1 vccd1 vccd1 _099_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_184_ _184_/A _102_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__ebufn_8
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_098_ _123_/A vssd1 vssd1 vccd1 vccd1 _103_/A sky130_fd_sc_hd__buf_6
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_167__66 vssd1 vssd1 vccd1 vccd1 _167__66/HI _200_/A sky130_fd_sc_hd__conb_1
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_137__36 vssd1 vssd1 vccd1 vccd1 _137__36/HI _170_/A sky130_fd_sc_hd__conb_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_183_ _183_/A _101_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__ebufn_8
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_151__50 vssd1 vssd1 vccd1 vccd1 _151__50/HI _184_/A sky130_fd_sc_hd__conb_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_097_ _097_/A vssd1 vssd1 vccd1 vccd1 _097_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_182_ _182_/A _100_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__ebufn_8
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_096_ _097_/A vssd1 vssd1 vccd1 vccd1 _096_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_158__57 vssd1 vssd1 vccd1 vccd1 _158__57/HI _191_/A sky130_fd_sc_hd__conb_1
XFILLER_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_181_ _181_/A _099_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__ebufn_8
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_142__41 vssd1 vssd1 vccd1 vccd1 _142__41/HI _175_/A sky130_fd_sc_hd__conb_1
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_095_ _097_/A vssd1 vssd1 vccd1 vccd1 _095_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_180_ _180_/A _097_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__ebufn_8
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_094_ _097_/A vssd1 vssd1 vccd1 vccd1 _094_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_129_ _129_/A _129_/B _129_/C _129_/D vssd1 vssd1 vccd1 vccd1 _135_/C sky130_fd_sc_hd__or4_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_149__48 vssd1 vssd1 vccd1 vccd1 _149__48/HI _182_/A sky130_fd_sc_hd__conb_1
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_163__62 vssd1 vssd1 vccd1 vccd1 _163__62/HI _196_/A sky130_fd_sc_hd__conb_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_093_ _097_/A vssd1 vssd1 vccd1 vccd1 _093_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput1 active vssd1 vssd1 vccd1 vccd1 _116_/A sky130_fd_sc_hd__buf_8
XFILLER_84_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_128_ _128_/A _128_/B _128_/C _128_/D vssd1 vssd1 vccd1 vccd1 _135_/B sky130_fd_sc_hd__or4_1
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_092_ _123_/A vssd1 vssd1 vccd1 vccd1 _097_/A sky130_fd_sc_hd__buf_4
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput2 wb_rst_i vssd1 vssd1 vccd1 vccd1 _124_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_127_ _127_/A _127_/B _127_/C vssd1 vssd1 vccd1 vccd1 _135_/A sky130_fd_sc_hd__or3_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_154__53 vssd1 vssd1 vccd1 vccd1 _154__53/HI _187_/A sky130_fd_sc_hd__conb_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_091_ _091_/A vssd1 vssd1 vccd1 vccd1 _091_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput3 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _129_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_126_ _126_/A _126_/B _126_/C _126_/D vssd1 vssd1 vccd1 vccd1 _127_/C sky130_fd_sc_hd__or4_4
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_109_ _109_/A vssd1 vssd1 vccd1 vccd1 _109_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_090_ _091_/A vssd1 vssd1 vccd1 vccd1 _090_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 _130_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_125_ _125_/A _125_/B input24/X input23/X vssd1 vssd1 vccd1 vccd1 _127_/B sky130_fd_sc_hd__or4bb_2
XFILLER_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_108_ _109_/A vssd1 vssd1 vccd1 vccd1 _108_/Y sky130_fd_sc_hd__inv_2
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_145__44 vssd1 vssd1 vccd1 vccd1 _145__44/HI _178_/A sky130_fd_sc_hd__conb_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput5 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 _131_/D sky130_fd_sc_hd__buf_4
XFILLER_110_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_124_ _124_/A _124_/B input35/X vssd1 vssd1 vccd1 vccd1 _127_/A sky130_fd_sc_hd__or3b_1
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput30 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _128_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_107_ _109_/A vssd1 vssd1 vccd1 vccd1 _107_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_160__59 vssd1 vssd1 vccd1 vccd1 _160__59/HI _193_/A sky130_fd_sc_hd__conb_1
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput6 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 _130_/C sky130_fd_sc_hd__buf_2
XFILLER_110_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_123_ _123_/A vssd1 vssd1 vccd1 vccd1 _123_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput20 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _126_/B sky130_fd_sc_hd__clkbuf_2
Xinput31 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _131_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_166__65 vssd1 vssd1 vccd1 vccd1 _166__65/HI _199_/A sky130_fd_sc_hd__conb_1
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_106_ _109_/A vssd1 vssd1 vccd1 vccd1 _106_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput7 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 _130_/B sky130_fd_sc_hd__buf_4
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_199_ _199_/A _120_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__ebufn_8
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_122_ _123_/A vssd1 vssd1 vccd1 vccd1 _122_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 _132_/C sky130_fd_sc_hd__buf_2
Xinput21 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _125_/A sky130_fd_sc_hd__clkbuf_4
Xinput32 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _128_/D sky130_fd_sc_hd__buf_2
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_105_ _109_/A vssd1 vssd1 vccd1 vccd1 _105_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 _132_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_198_ _198_/A _119_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__ebufn_8
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_121_ _121_/A vssd1 vssd1 vccd1 vccd1 _121_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _126_/D sky130_fd_sc_hd__buf_2
Xinput11 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _132_/B sky130_fd_sc_hd__clkbuf_4
Xinput33 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _131_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_104_ _116_/A vssd1 vssd1 vccd1 vccd1 _109_/A sky130_fd_sc_hd__buf_6
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_157__56 vssd1 vssd1 vccd1 vccd1 _157__56/HI _190_/A sky130_fd_sc_hd__conb_1
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_141__40 vssd1 vssd1 vccd1 vccd1 _141__40/HI _174_/A sky130_fd_sc_hd__conb_1
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _130_/D sky130_fd_sc_hd__buf_4
XFILLER_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_197_ _197_/A _118_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__ebufn_8
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_120_ _121_/A vssd1 vssd1 vccd1 vccd1 _120_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _133_/A sky130_fd_sc_hd__buf_2
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput34 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _131_/B sky130_fd_sc_hd__clkbuf_4
Xinput23 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_2
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_103_ _103_/A vssd1 vssd1 vccd1 vccd1 _103_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_196_ _196_/A _117_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__ebufn_8
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _132_/D sky130_fd_sc_hd__buf_2
Xinput35 wbs_stb_i vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_4
Xinput24 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_179_ _179_/A _096_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__ebufn_8
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_102_ _103_/A vssd1 vssd1 vccd1 vccd1 _102_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_148__47 vssd1 vssd1 vccd1 vccd1 _148__47/HI _181_/A sky130_fd_sc_hd__conb_1
XFILLER_92_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_162__61 vssd1 vssd1 vccd1 vccd1 _162__61/HI _195_/A sky130_fd_sc_hd__conb_1
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_195_ _195_/A _115_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__ebufn_8
XFILLER_123_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput14 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _129_/B sky130_fd_sc_hd__buf_4
Xinput25 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _128_/A sky130_fd_sc_hd__clkbuf_4
X_178_ _178_/A _095_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__ebufn_8
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_101_ _103_/A vssd1 vssd1 vccd1 vccd1 _101_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_194_ _194_/A _114_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__ebufn_8
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput26 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 _124_/A sky130_fd_sc_hd__clkbuf_2
Xinput15 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _133_/C sky130_fd_sc_hd__buf_2
X_177_ _177_/A _094_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__ebufn_8
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_100_ _103_/A vssd1 vssd1 vccd1 vccd1 _100_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_139__38 vssd1 vssd1 vccd1 vccd1 _139__38/HI _172_/A sky130_fd_sc_hd__conb_1
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_153__52 vssd1 vssd1 vccd1 vccd1 _153__52/HI _186_/A sky130_fd_sc_hd__conb_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_193_ _193_/A _113_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__ebufn_8
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _133_/B sky130_fd_sc_hd__clkbuf_4
Xinput27 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 _125_/B sky130_fd_sc_hd__buf_2
X_176_ _176_/A _093_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__ebufn_8
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_192_ _192_/A _112_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__ebufn_8
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput28 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _129_/D sky130_fd_sc_hd__buf_2
Xinput17 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 _126_/A sky130_fd_sc_hd__buf_2
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_175_ _175_/A _091_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__ebufn_8
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_089_ _091_/A vssd1 vssd1 vccd1 vccd1 _089_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_144__43 vssd1 vssd1 vccd1 vccd1 _144__43/HI _177_/A sky130_fd_sc_hd__conb_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_191_ _191_/A _111_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__ebufn_8
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput18 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _133_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput29 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _128_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_174_ _174_/A _090_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__ebufn_8
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_088_ _091_/A vssd1 vssd1 vccd1 vccd1 _088_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_190_ _190_/A _109_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__ebufn_8
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput19 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _126_/C sky130_fd_sc_hd__clkbuf_2
X_173_ _173_/A _089_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__ebufn_8
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_165__64 vssd1 vssd1 vccd1 vccd1 _165__64/HI _198_/A sky130_fd_sc_hd__conb_1
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_087_ _091_/A vssd1 vssd1 vccd1 vccd1 _087_/Y sky130_fd_sc_hd__inv_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_172_ _172_/A _088_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__ebufn_8
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_086_ _123_/A vssd1 vssd1 vccd1 vccd1 _091_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_150__49 vssd1 vssd1 vccd1 vccd1 _150__49/HI _183_/A sky130_fd_sc_hd__conb_1
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_171_ _171_/A _087_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__ebufn_8
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_085_ _116_/A vssd1 vssd1 vccd1 vccd1 _123_/A sky130_fd_sc_hd__buf_6
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_156__55 vssd1 vssd1 vccd1 vccd1 _156__55/HI _189_/A sky130_fd_sc_hd__conb_1
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_170_ _170_/A _123_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__ebufn_8
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_084_ _116_/A vssd1 vssd1 vccd1 vccd1 _129_/A sky130_fd_sc_hd__inv_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_136_ wb_clk_i _136_/D vssd1 vssd1 vccd1 vccd1 _169_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_119_ _121_/A vssd1 vssd1 vccd1 vccd1 _119_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_0 wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_147__46 vssd1 vssd1 vccd1 vccd1 _147__46/HI _180_/A sky130_fd_sc_hd__conb_1
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_161__60 vssd1 vssd1 vccd1 vccd1 _161__60/HI _194_/A sky130_fd_sc_hd__conb_1
X_135_ _135_/A _135_/B _135_/C _135_/D vssd1 vssd1 vccd1 vccd1 _136_/D sky130_fd_sc_hd__nor4_1
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_118_ _121_/A vssd1 vssd1 vccd1 vccd1 _118_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_1 wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_134_ _134_/A _134_/B _134_/C _134_/D vssd1 vssd1 vccd1 vccd1 _135_/D sky130_fd_sc_hd__or4_1
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_117_ _121_/A vssd1 vssd1 vccd1 vccd1 _117_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_2 _133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_168__67 vssd1 vssd1 vccd1 vccd1 _168__67/HI _201_/A sky130_fd_sc_hd__conb_1
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_138__37 vssd1 vssd1 vccd1 vccd1 _138__37/HI _171_/A sky130_fd_sc_hd__conb_1
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_133_ _133_/A _133_/B _133_/C _133_/D vssd1 vssd1 vccd1 vccd1 _134_/D sky130_fd_sc_hd__or4_1
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_152__51 vssd1 vssd1 vccd1 vccd1 _152__51/HI _185_/A sky130_fd_sc_hd__conb_1
XFILLER_115_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_116_ _116_/A vssd1 vssd1 vccd1 vccd1 _121_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_3 _125_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_201_ _201_/A _122_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__ebufn_8
X_132_ _132_/A _132_/B _132_/C _132_/D vssd1 vssd1 vccd1 vccd1 _134_/C sky130_fd_sc_hd__or4_1
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_115_ _115_/A vssd1 vssd1 vccd1 vccd1 _115_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
.ends

